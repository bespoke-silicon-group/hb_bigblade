
module bsg_chip_core_complex

 import bsg_chip_pkg::*;
 import bsg_noc_pkg::*;
 import bsg_manycore_pkg::*;

  (input                      hb_clk_i
  ,input                      router_clk_i
  ,input bsg_chip_tag_lines_s tag_lines_i

  ,input  bsg_chip_io_link_sif_s [io_link_num_gp-1:0][io_ct_num_in_gp-1:0] io_links_i
  ,output bsg_chip_io_link_sif_s [io_link_num_gp-1:0][io_ct_num_in_gp-1:0] io_links_o

  ,input  bsg_chip_mem_link_sif_s [mem_link_num_gp-1:0] mem_links_i
  ,output bsg_chip_mem_link_sif_s [mem_link_num_gp-1:0] mem_links_o
  );

  //////////////////////////////////////////////////
  //
  // BSG Tag Client Instance
  //

  // Tag payload for hb control signals
  typedef struct packed { 
      logic padding;
      logic reset;
  } hb_tag_payload_s;

  hb_tag_payload_s hb_tag_data_lo;
  logic            hb_tag_new_data_lo;

  bsg_tag_client #(.width_p( $bits(hb_tag_data_lo) ), .default_p( 0 ))
    btc_hb
      (.bsg_tag_i     ( tag_lines_i.hb_reset )
      ,.recv_clk_i    ( hb_clk_i )
      ,.recv_reset_i  ( 1'b0 )
      ,.recv_new_r_o  ( hb_tag_new_data_lo )
      ,.recv_data_r_o ( hb_tag_data_lo )
      );

  // Tag payload for router control signals
  typedef struct packed { 
      logic padding;
      logic reset;
  } router_tag_payload_s;

  router_tag_payload_s router_tag_data_lo;
  logic                router_tag_new_data_lo;

  bsg_tag_client #(.width_p( $bits(router_tag_data_lo) ), .default_p( 0 ))
    btc_router
      (.bsg_tag_i     ( tag_lines_i.router_reset )
      ,.recv_clk_i    ( router_clk_i )
      ,.recv_reset_i  ( 1'b0 )
      ,.recv_new_r_o  ( router_tag_new_data_lo )
      ,.recv_data_r_o ( router_tag_data_lo )
      );


  //////////////////////////////////////////////////
  //
  // Manycore Array
  //
  `declare_bsg_manycore_link_sif_s(hb_addr_width_gp,hb_data_width_gp,hb_x_cord_width_gp,hb_y_cord_width_gp);
  `declare_bsg_manycore_ruche_x_link_sif_s(hb_addr_width_gp,hb_data_width_gp,hb_x_cord_width_gp,hb_y_cord_width_gp);
  `declare_bsg_ready_and_link_sif_s(wh_flit_width_gp, wh_link_sif_s);

  bsg_manycore_link_sif_s [(hb_num_pods_x_gp*hb_num_tiles_x_gp)-1:0] io_link_sif_li;
  bsg_manycore_link_sif_s [(hb_num_pods_x_gp*hb_num_tiles_x_gp)-1:0] io_link_sif_lo;
  wh_link_sif_s [E:W][hb_num_pods_y_gp-1:0][S:N][wh_ruche_factor_gp-1:0] wh_unconc_link_sif_li;
  wh_link_sif_s [E:W][hb_num_pods_y_gp-1:0][S:N][wh_ruche_factor_gp-1:0] wh_unconc_link_sif_lo;
  bsg_manycore_link_sif_s [E:W][hb_num_pods_y_gp-1:0][hb_num_tiles_y_gp-1:0] hor_link_sif_li;
  bsg_manycore_link_sif_s [E:W][hb_num_pods_y_gp-1:0][hb_num_tiles_y_gp-1:0] hor_link_sif_lo;
  bsg_manycore_ruche_x_link_sif_s [E:W][hb_num_pods_y_gp-1:0][hb_num_tiles_y_gp-1:0][hb_ruche_factor_X_gp-1:0] ruche_link_li;
  bsg_manycore_ruche_x_link_sif_s [E:W][hb_num_pods_y_gp-1:0][hb_num_tiles_y_gp-1:0][hb_ruche_factor_X_gp-1:0] ruche_link_lo;

  bsg_manycore_pod_ruche_array #(
    .num_tiles_x_p(hb_num_tiles_x_gp)
    ,.num_tiles_y_p(hb_num_tiles_y_gp)
    ,.pod_x_cord_width_p(hb_pod_x_cord_width_gp)
    ,.pod_y_cord_width_p(hb_pod_y_cord_width_gp)
    ,.x_cord_width_p(hb_x_cord_width_gp)
    ,.y_cord_width_p(hb_y_cord_width_gp)
    ,.addr_width_p(hb_addr_width_gp)
    ,.data_width_p(hb_data_width_gp)
    ,.ruche_factor_X_p(hb_ruche_factor_X_gp)
    
    ,.dmem_size_p(hb_dmem_size_gp)
    ,.icache_entries_p(hb_icache_entries_gp)
    ,.icache_tag_width_p(hb_icache_tag_width_gp)

    ,.vcache_addr_width_p(vcache_addr_width_gp)
    ,.vcache_data_width_p(vcache_data_width_gp)
    ,.vcache_ways_p(vcache_ways_gp)
    ,.vcache_sets_p(vcache_sets_gp)
    ,.vcache_block_size_in_words_p(vcache_block_size_in_words_gp)
    ,.vcache_size_p(vcache_size_gp)
    ,.vcache_dma_data_width_p(vcache_dma_data_width_gp)

    ,.wh_ruche_factor_p(wh_ruche_factor_gp)
    ,.wh_cid_width_p(wh_cid_width_gp)
    ,.wh_flit_width_p(wh_flit_width_gp)
    ,.wh_cord_width_p(wh_cord_width_gp)
    ,.wh_len_width_p(wh_len_width_gp)

    ,.num_pods_y_p(hb_num_pods_y_gp)
    ,.num_pods_x_p(hb_num_pods_x_gp)

    ,.reset_depth_p(hb_reset_depth_gp)
  ) DUT (
    .clk_i(hb_clk_i)
    ,.reset_i(hb_tag_data_lo.reset)

    ,.io_link_sif_i(io_link_sif_li)
    ,.io_link_sif_o(io_link_sif_lo)

    ,.wh_link_sif_i(wh_unconc_link_sif_li)
    ,.wh_link_sif_o(wh_unconc_link_sif_lo)

    ,.hor_link_sif_i(hor_link_sif_li)
    ,.hor_link_sif_o(hor_link_sif_lo)

    ,.ruche_link_i(ruche_link_li)
    ,.ruche_link_o(ruche_link_lo)

    ,.bsg_tag_i(tag_lines_i.hb_pod)
  );

  // hor tieoff
  for (genvar i = W; i <= E; i++) begin
    for (genvar j = 0; j < hb_num_pods_y_gp; j++) begin
      for (genvar k = 0; k < hb_num_tiles_y_gp; k++) begin
        bsg_manycore_link_sif_tieoff #(
          .addr_width_p(hb_addr_width_gp)
          ,.data_width_p(hb_data_width_gp)
          ,.x_cord_width_p(hb_x_cord_width_gp)
          ,.y_cord_width_p(hb_y_cord_width_gp)
        ) hor_tieoff (
          .clk_i(hb_clk_i)
          ,.reset_i(hb_tag_data_lo.reset)
          ,.link_sif_i(hor_link_sif_lo[i][j][k])
          ,.link_sif_o(hor_link_sif_li[i][j][k])
        );
      end
    end
  end

  // ruche tieoff
  for (genvar i = W; i <= E; i++) begin
    for (genvar j = 0; j < hb_num_pods_y_gp; j++) begin
      for (genvar k = 0; k < hb_num_tiles_y_gp; k++) begin
        for (genvar l = 0; l < hb_ruche_factor_X_gp; l++) begin
          bsg_manycore_ruche_x_link_sif_tieoff #(
            .addr_width_p(hb_addr_width_gp)
            ,.data_width_p(hb_data_width_gp)
            ,.x_cord_width_p(hb_x_cord_width_gp)
            ,.y_cord_width_p(hb_y_cord_width_gp)
            ,.ruche_stage_p(l)
            ,.ruche_factor_X_p(hb_ruche_factor_X_gp)
            ,.west_not_east_p(i==W ? 1 : 0)
          ) ruche_tieoff (
            .clk_i(hb_clk_i)
            ,.reset_i(hb_tag_data_lo.reset)
            ,.ruche_link_i(ruche_link_lo[i][j][k][l])
            ,.ruche_link_o(ruche_link_li[i][j][k][l]) 
          );
        end  
      end
    end
  end


  // io tieoff
  for (genvar i = 1; i < hb_num_pods_x_gp*hb_num_tiles_x_gp; i++) begin
    bsg_manycore_link_sif_tieoff #(
      .addr_width_p(hb_addr_width_gp)
      ,.data_width_p(hb_data_width_gp)
      ,.x_cord_width_p(hb_x_cord_width_gp)
      ,.y_cord_width_p(hb_y_cord_width_gp)
    ) io_n_tieoff (
      .clk_i(hb_clk_i)
      ,.reset_i(hb_tag_data_lo.reset)
      ,.link_sif_i(io_link_sif_lo[i])
      ,.link_sif_o(io_link_sif_li[i])
    );
  end


  //////////////////////////////////////////////////
  //
  // Manycore Adapter
  //
  bsg_manycore_link_sif_s [io_link_num_gp-1:0] manycore_links_li;
  bsg_manycore_link_sif_s [io_link_num_gp-1:0] manycore_links_lo;
  
  assign io_link_sif_li[0] = manycore_links_li[0];
  assign manycore_links_lo = {'0, io_link_sif_lo[0]};
  
  for (genvar i = 0; i < io_link_num_gp; i++)
  begin: mc_io
    bsg_manycore_link_async_to_bsg_link
   #(.addr_width_p    (hb_addr_width_gp  )
    ,.data_width_p    (hb_data_width_gp  )
    ,.x_cord_width_p  (hb_x_cord_width_gp)
    ,.y_cord_width_p  (hb_y_cord_width_gp)
    ,.bsg_link_width_p(io_ct_width_gp    )
    ) mc_adapter
    (.mc_clk_i        (hb_clk_i)
    ,.mc_reset_i      (hb_tag_data_lo.reset)
    ,.mc_links_sif_i  (manycore_links_lo[i])
    ,.mc_links_sif_o  (manycore_links_li[i])
  
    ,.bsg_link_clk_i  (router_clk_i)
    ,.bsg_link_reset_i(router_tag_data_lo.reset)
    ,.bsg_link_i      (io_links_i[i])
    ,.bsg_link_o      (io_links_o[i])
    );
  end


  // clock domain crossing
  wh_link_sif_s [E:W][hb_num_pods_y_gp-1:0][S:N][wh_ruche_factor_gp-1:0] router_unconc_link_sif_li;
  wh_link_sif_s [E:W][hb_num_pods_y_gp-1:0][S:N][wh_ruche_factor_gp-1:0] router_unconc_link_sif_lo;
  for (genvar i = W; i <= E; i++) begin: cdc_s
    for (genvar j = 0; j < hb_num_pods_y_gp; j++) begin: cdc_y
      for (genvar m = N; m <= S; m++) begin: cdc_tb
        for (genvar l = 0; l < wh_ruche_factor_gp; l++) begin: cdc_f
          bsg_ready_and_link_async_to_bsg_link
         #(.ral_link_width_p(wh_flit_width_gp)
          ,.bsg_link_width_p(wh_flit_width_gp)
          ) async
          (.ral_clk_i       (hb_clk_i)
          ,.ral_reset_i     (hb_tag_data_lo.reset)
          ,.ral_link_i      (wh_unconc_link_sif_lo[i][j][m][l])
          ,.ral_link_o      (wh_unconc_link_sif_li[i][j][m][l])
          ,.bsg_link_clk_i  (router_clk_i)
          ,.bsg_link_reset_i(router_tag_data_lo.reset)
          ,.bsg_link_i      (router_unconc_link_sif_li[i][j][m][l])
          ,.bsg_link_o      (router_unconc_link_sif_lo[i][j][m][l])
          );
        end
      end
    end
  end

  // instantiate wormhole concentrators
  wh_link_sif_s [E:W][hb_num_pods_y_gp-1:0] wh_link_sif_li;
  wh_link_sif_s [E:W][hb_num_pods_y_gp-1:0] wh_link_sif_lo;

  for (genvar i = W; i <= E; i++) begin: conc_s
    for (genvar j = 0; j < hb_num_pods_y_gp; j++) begin: conc_y
      bsg_wormhole_concentrator #(
        .flit_width_p(wh_flit_width_gp)
        ,.len_width_p(wh_len_width_gp)
        ,.cid_width_p(wh_cid_width_gp)
        ,.cord_width_p(wh_cord_width_gp)
        ,.num_in_p(2*wh_ruche_factor_gp)
      ) conc0 (
        .clk_i(router_clk_i)
        ,.reset_i(router_tag_data_lo.reset)
      
        ,.links_i(router_unconc_link_sif_lo[i][j])
        ,.links_o(router_unconc_link_sif_li[i][j])

        ,.concentrated_link_i(wh_link_sif_li[i][j])
        ,.concentrated_link_o(wh_link_sif_lo[i][j])
      );
    end
  end

  // Attach wormhole links to mem links
  bsg_chip_mem_link_sif_s [mem_link_conc_num_gp-1:0] mem_links_conc_li;
  bsg_chip_mem_link_sif_s [mem_link_conc_num_gp-1:0] mem_links_conc_lo;

  for (genvar i = 0; i < mem_link_conc_num_gp/2; i++) begin
    if (i < hb_num_pods_y_gp) begin
      assign wh_link_sif_li[W][i].v             = mem_links_conc_li[i].v;
      assign wh_link_sif_li[W][i].data          = mem_links_conc_li[i].data;
      assign wh_link_sif_li[W][i].ready_and_rev = mem_links_conc_li[i].ready_and_rev;
      assign mem_links_conc_lo[i].v             = wh_link_sif_lo[W][i].v;
      assign mem_links_conc_lo[i].data          = wh_link_sif_lo[W][i].data;
      assign mem_links_conc_lo[i].ready_and_rev = wh_link_sif_lo[W][i].ready_and_rev;
      assign wh_link_sif_li[E][i].v             = mem_links_conc_li[i+mem_link_conc_num_gp/2].v;
      assign wh_link_sif_li[E][i].data          = mem_links_conc_li[i+mem_link_conc_num_gp/2].data;
      assign wh_link_sif_li[E][i].ready_and_rev = mem_links_conc_li[i+mem_link_conc_num_gp/2].ready_and_rev;
      assign mem_links_conc_lo[i+mem_link_conc_num_gp/2].v             = wh_link_sif_lo[E][i].v;
      assign mem_links_conc_lo[i+mem_link_conc_num_gp/2].data          = wh_link_sif_lo[E][i].data;
      assign mem_links_conc_lo[i+mem_link_conc_num_gp/2].ready_and_rev = wh_link_sif_lo[E][i].ready_and_rev;
    end else begin
      assign mem_links_conc_lo[i] = '0;
      assign mem_links_conc_lo[i+mem_link_conc_num_gp/2] = '0;
    end
  end

  // mem link round robin arbiters
  for (genvar i = 0; i < mem_link_conc_num_gp; i++) begin: mem_link_arb
    bsg_ready_and_link_round_robin_static 
   #(.width_p      (mem_link_width_gp   )
    ,.num_in_p     (mem_link_rr_ratio_gp)
    ) rr
    (.clk_i        (router_clk_i        )
    ,.reset_i      (router_tag_data_lo.reset)
    ,.single_link_i(mem_links_conc_lo[i])
    ,.single_link_o(mem_links_conc_li[i])
    ,.links_i      (mem_links_i[i*mem_link_rr_ratio_gp+:mem_link_rr_ratio_gp])
    ,.links_o      (mem_links_o[i*mem_link_rr_ratio_gp+:mem_link_rr_ratio_gp])
    );
  end

endmodule