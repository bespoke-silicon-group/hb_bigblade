// bsg_hb_pcb.v
//
// simulates connectivity of the asic cloud PCB
//
// this is intended as the canonical simulation file
// but currently it may only implement a subset of
// all of the wires and functionality -- please
// extend rather than cloning the file and modifying it
//

`timescale 1ps/1ps

module bsg_hb_pcb
(
    // this is the FMC connector
    inout [33:00] LAxx_N
    , inout [33:00] LAxx_P      //  e.g. LA14_N
    , inout CLK0_C2M_N
    , inout CLK0_C2M_P
    , inout CLK0_M2C_N
    , inout CLK0_M2C_P

    // SMA connectors (for simulation)
    , input ASIC_SMA_IN_N
    , input ASIC_SMA_IN_P       // terminated on ASIC side
    , inout ASIC_SMA_OUT_N
    , inout ASIC_SMA_OUT_P      // unterminated

    , inout FPGA_SMA_IN_N
    , inout FPGA_SMA_IN_P       // unterminated
    , inout FPGA_SMA_OUT_N
    , inout FPGA_SMA_OUT_P      // unterminated

    // LEDs (for simulation)
    , output [3:0] FPGA_LED     // from GW   FPGA
    , output [1:0] ASIC_LED     // from ASIC FPGA

    , input  UART_RX
    , output UART_TX

    // low-true reset signal for GW FPGA (normal driven by reset controller)
    , input PWR_RSTN
  );


  //
  // Comm link wires (Between GW and IC)
  //

  wire [19:0] IC_GW_LINK_CLK;
  wire [19:0] IC_GW_LINK_V;
  wire [19:0] IC_GW_LINK_TKN;
  wire [19:0] IC_GW_LINK_D0;
  wire [19:0] IC_GW_LINK_D1;
  wire [19:0] IC_GW_LINK_D2;
  wire [19:0] IC_GW_LINK_D3;
  wire [19:0] IC_GW_LINK_D4;
  wire [19:0] IC_GW_LINK_D5;
  wire [19:0] IC_GW_LINK_D6;
  wire [19:0] IC_GW_LINK_D7;
  wire [19:0] IC_GW_LINK_D8;

  wire [19:0] GW_IC_LINK_CLK;
  wire [19:0] GW_IC_LINK_V;
  wire [19:0] GW_IC_LINK_TKN;
  wire [19:0] GW_IC_LINK_D0;
  wire [19:0] GW_IC_LINK_D1;
  wire [19:0] GW_IC_LINK_D2;
  wire [19:0] GW_IC_LINK_D3;
  wire [19:0] GW_IC_LINK_D4;
  wire [19:0] GW_IC_LINK_D5;
  wire [19:0] GW_IC_LINK_D6;
  wire [19:0] GW_IC_LINK_D7;
  wire [19:0] GW_IC_LINK_D8;


  //
  // Misc wires (GW)
  //
  wire GW_TAG_CLKO;
  wire GW_TAG_DATAO;
  wire GW_TAG_EN;

  wire GW_CLKA;
  wire GW_CLKB;
  wire GW_CLKC;

  wire GW_SEL0;
  wire GW_SEL1;
  //wire GW_SEL2;

  wire GW_CLK_RESET;
  wire GW_CORE_RESET;


  //
  // Misc wires (IC)
  //
  wire IC_CLKO;  // Clock out (for scoping clock generators)

  //
  // GATEWAY SOCKET
  //

  bsg_gateway_chip GW
  (.p_bsg_link_in0_clk_o (GW_IC_LINK_CLK  [0])
  ,.p_bsg_link_in0_v_o   (GW_IC_LINK_V    [0])
  ,.p_bsg_link_in0_tkn_i (GW_IC_LINK_TKN  [0])
  ,.p_bsg_link_in0_d0_o  (GW_IC_LINK_D0   [0])
  ,.p_bsg_link_in0_d1_o  (GW_IC_LINK_D1   [0])
  ,.p_bsg_link_in0_d2_o  (GW_IC_LINK_D2   [0])
  ,.p_bsg_link_in0_d3_o  (GW_IC_LINK_D3   [0])
  ,.p_bsg_link_in0_d4_o  (GW_IC_LINK_D4   [0])
  ,.p_bsg_link_in0_d5_o  (GW_IC_LINK_D5   [0])
  ,.p_bsg_link_in0_d6_o  (GW_IC_LINK_D6   [0])
  ,.p_bsg_link_in0_d7_o  (GW_IC_LINK_D7   [0])
  ,.p_bsg_link_in0_d8_o  (GW_IC_LINK_D8   [0])
                          
  ,.p_bsg_link_in1_clk_o (GW_IC_LINK_CLK  [1])
  ,.p_bsg_link_in1_v_o   (GW_IC_LINK_V    [1])
  ,.p_bsg_link_in1_tkn_i (GW_IC_LINK_TKN  [1])
  ,.p_bsg_link_in1_d0_o  (GW_IC_LINK_D0   [1])
  ,.p_bsg_link_in1_d1_o  (GW_IC_LINK_D1   [1])
  ,.p_bsg_link_in1_d2_o  (GW_IC_LINK_D2   [1])
  ,.p_bsg_link_in1_d3_o  (GW_IC_LINK_D3   [1])
  ,.p_bsg_link_in1_d4_o  (GW_IC_LINK_D4   [1])
  ,.p_bsg_link_in1_d5_o  (GW_IC_LINK_D5   [1])
  ,.p_bsg_link_in1_d6_o  (GW_IC_LINK_D6   [1])
  ,.p_bsg_link_in1_d7_o  (GW_IC_LINK_D7   [1])
  ,.p_bsg_link_in1_d8_o  (GW_IC_LINK_D8   [1])
                          
  ,.p_bsg_link_in2_clk_o (GW_IC_LINK_CLK  [2])
  ,.p_bsg_link_in2_v_o   (GW_IC_LINK_V    [2])
  ,.p_bsg_link_in2_tkn_i (GW_IC_LINK_TKN  [2])
  ,.p_bsg_link_in2_d0_o  (GW_IC_LINK_D0   [2])
  ,.p_bsg_link_in2_d1_o  (GW_IC_LINK_D1   [2])
  ,.p_bsg_link_in2_d2_o  (GW_IC_LINK_D2   [2])
  ,.p_bsg_link_in2_d3_o  (GW_IC_LINK_D3   [2])
  ,.p_bsg_link_in2_d4_o  (GW_IC_LINK_D4   [2])
  ,.p_bsg_link_in2_d5_o  (GW_IC_LINK_D5   [2])
  ,.p_bsg_link_in2_d6_o  (GW_IC_LINK_D6   [2])
  ,.p_bsg_link_in2_d7_o  (GW_IC_LINK_D7   [2])
  ,.p_bsg_link_in2_d8_o  (GW_IC_LINK_D8   [2])
                          
  ,.p_bsg_link_in3_clk_o (GW_IC_LINK_CLK  [3])
  ,.p_bsg_link_in3_v_o   (GW_IC_LINK_V    [3])
  ,.p_bsg_link_in3_tkn_i (GW_IC_LINK_TKN  [3])
  ,.p_bsg_link_in3_d0_o  (GW_IC_LINK_D0   [3])
  ,.p_bsg_link_in3_d1_o  (GW_IC_LINK_D1   [3])
  ,.p_bsg_link_in3_d2_o  (GW_IC_LINK_D2   [3])
  ,.p_bsg_link_in3_d3_o  (GW_IC_LINK_D3   [3])
  ,.p_bsg_link_in3_d4_o  (GW_IC_LINK_D4   [3])
  ,.p_bsg_link_in3_d5_o  (GW_IC_LINK_D5   [3])
  ,.p_bsg_link_in3_d6_o  (GW_IC_LINK_D6   [3])
  ,.p_bsg_link_in3_d7_o  (GW_IC_LINK_D7   [3])
  ,.p_bsg_link_in3_d8_o  (GW_IC_LINK_D8   [3])
                          
  ,.p_bsg_link_in4_clk_o (GW_IC_LINK_CLK  [4])
  ,.p_bsg_link_in4_v_o   (GW_IC_LINK_V    [4])
  ,.p_bsg_link_in4_tkn_i (GW_IC_LINK_TKN  [4])
  ,.p_bsg_link_in4_d0_o  (GW_IC_LINK_D0   [4])
  ,.p_bsg_link_in4_d1_o  (GW_IC_LINK_D1   [4])
  ,.p_bsg_link_in4_d2_o  (GW_IC_LINK_D2   [4])
  ,.p_bsg_link_in4_d3_o  (GW_IC_LINK_D3   [4])
  ,.p_bsg_link_in4_d4_o  (GW_IC_LINK_D4   [4])
  ,.p_bsg_link_in4_d5_o  (GW_IC_LINK_D5   [4])
  ,.p_bsg_link_in4_d6_o  (GW_IC_LINK_D6   [4])
  ,.p_bsg_link_in4_d7_o  (GW_IC_LINK_D7   [4])
  ,.p_bsg_link_in4_d8_o  (GW_IC_LINK_D8   [4])
                          
  ,.p_bsg_link_in5_clk_o (GW_IC_LINK_CLK  [5])
  ,.p_bsg_link_in5_v_o   (GW_IC_LINK_V    [5])
  ,.p_bsg_link_in5_tkn_i (GW_IC_LINK_TKN  [5])
  ,.p_bsg_link_in5_d0_o  (GW_IC_LINK_D0   [5])
  ,.p_bsg_link_in5_d1_o  (GW_IC_LINK_D1   [5])
  ,.p_bsg_link_in5_d2_o  (GW_IC_LINK_D2   [5])
  ,.p_bsg_link_in5_d3_o  (GW_IC_LINK_D3   [5])
  ,.p_bsg_link_in5_d4_o  (GW_IC_LINK_D4   [5])
  ,.p_bsg_link_in5_d5_o  (GW_IC_LINK_D5   [5])
  ,.p_bsg_link_in5_d6_o  (GW_IC_LINK_D6   [5])
  ,.p_bsg_link_in5_d7_o  (GW_IC_LINK_D7   [5])
  ,.p_bsg_link_in5_d8_o  (GW_IC_LINK_D8   [5])
                           
  ,.p_bsg_link_in6_clk_o (GW_IC_LINK_CLK  [6])
  ,.p_bsg_link_in6_v_o   (GW_IC_LINK_V    [6])
  ,.p_bsg_link_in6_tkn_i (GW_IC_LINK_TKN  [6])
  ,.p_bsg_link_in6_d0_o  (GW_IC_LINK_D0   [6])
  ,.p_bsg_link_in6_d1_o  (GW_IC_LINK_D1   [6])
  ,.p_bsg_link_in6_d2_o  (GW_IC_LINK_D2   [6])
  ,.p_bsg_link_in6_d3_o  (GW_IC_LINK_D3   [6])
  ,.p_bsg_link_in6_d4_o  (GW_IC_LINK_D4   [6])
  ,.p_bsg_link_in6_d5_o  (GW_IC_LINK_D5   [6])
  ,.p_bsg_link_in6_d6_o  (GW_IC_LINK_D6   [6])
  ,.p_bsg_link_in6_d7_o  (GW_IC_LINK_D7   [6])
  ,.p_bsg_link_in6_d8_o  (GW_IC_LINK_D8   [6])
                           
  ,.p_bsg_link_in7_clk_o (GW_IC_LINK_CLK  [7])
  ,.p_bsg_link_in7_v_o   (GW_IC_LINK_V    [7])
  ,.p_bsg_link_in7_tkn_i (GW_IC_LINK_TKN  [7])
  ,.p_bsg_link_in7_d0_o  (GW_IC_LINK_D0   [7])
  ,.p_bsg_link_in7_d1_o  (GW_IC_LINK_D1   [7])
  ,.p_bsg_link_in7_d2_o  (GW_IC_LINK_D2   [7])
  ,.p_bsg_link_in7_d3_o  (GW_IC_LINK_D3   [7])
  ,.p_bsg_link_in7_d4_o  (GW_IC_LINK_D4   [7])
  ,.p_bsg_link_in7_d5_o  (GW_IC_LINK_D5   [7])
  ,.p_bsg_link_in7_d6_o  (GW_IC_LINK_D6   [7])
  ,.p_bsg_link_in7_d7_o  (GW_IC_LINK_D7   [7])
  ,.p_bsg_link_in7_d8_o  (GW_IC_LINK_D8   [7])
                           
  ,.p_bsg_link_in8_clk_o (GW_IC_LINK_CLK  [8])
  ,.p_bsg_link_in8_v_o   (GW_IC_LINK_V    [8])
  ,.p_bsg_link_in8_tkn_i (GW_IC_LINK_TKN  [8])
  ,.p_bsg_link_in8_d0_o  (GW_IC_LINK_D0   [8])
  ,.p_bsg_link_in8_d1_o  (GW_IC_LINK_D1   [8])
  ,.p_bsg_link_in8_d2_o  (GW_IC_LINK_D2   [8])
  ,.p_bsg_link_in8_d3_o  (GW_IC_LINK_D3   [8])
  ,.p_bsg_link_in8_d4_o  (GW_IC_LINK_D4   [8])
  ,.p_bsg_link_in8_d5_o  (GW_IC_LINK_D5   [8])
  ,.p_bsg_link_in8_d6_o  (GW_IC_LINK_D6   [8])
  ,.p_bsg_link_in8_d7_o  (GW_IC_LINK_D7   [8])
  ,.p_bsg_link_in8_d8_o  (GW_IC_LINK_D8   [8])
                           
  ,.p_bsg_link_in9_clk_o (GW_IC_LINK_CLK  [9])
  ,.p_bsg_link_in9_v_o   (GW_IC_LINK_V    [9])
  ,.p_bsg_link_in9_tkn_i (GW_IC_LINK_TKN  [9])
  ,.p_bsg_link_in9_d0_o  (GW_IC_LINK_D0   [9])
  ,.p_bsg_link_in9_d1_o  (GW_IC_LINK_D1   [9])
  ,.p_bsg_link_in9_d2_o  (GW_IC_LINK_D2   [9])
  ,.p_bsg_link_in9_d3_o  (GW_IC_LINK_D3   [9])
  ,.p_bsg_link_in9_d4_o  (GW_IC_LINK_D4   [9])
  ,.p_bsg_link_in9_d5_o  (GW_IC_LINK_D5   [9])
  ,.p_bsg_link_in9_d6_o  (GW_IC_LINK_D6   [9])
  ,.p_bsg_link_in9_d7_o  (GW_IC_LINK_D7   [9])
  ,.p_bsg_link_in9_d8_o  (GW_IC_LINK_D8   [9])
                          
  ,.p_bsg_link_in10_clk_o(GW_IC_LINK_CLK  [10])
  ,.p_bsg_link_in10_v_o  (GW_IC_LINK_V    [10])
  ,.p_bsg_link_in10_tkn_i(GW_IC_LINK_TKN  [10])
  ,.p_bsg_link_in10_d0_o (GW_IC_LINK_D0   [10])
  ,.p_bsg_link_in10_d1_o (GW_IC_LINK_D1   [10])
  ,.p_bsg_link_in10_d2_o (GW_IC_LINK_D2   [10])
  ,.p_bsg_link_in10_d3_o (GW_IC_LINK_D3   [10])
  ,.p_bsg_link_in10_d4_o (GW_IC_LINK_D4   [10])
  ,.p_bsg_link_in10_d5_o (GW_IC_LINK_D5   [10])
  ,.p_bsg_link_in10_d6_o (GW_IC_LINK_D6   [10])
  ,.p_bsg_link_in10_d7_o (GW_IC_LINK_D7   [10])
  ,.p_bsg_link_in10_d8_o (GW_IC_LINK_D8   [10])
                           
  ,.p_bsg_link_in11_clk_o(GW_IC_LINK_CLK  [11])
  ,.p_bsg_link_in11_v_o  (GW_IC_LINK_V    [11])
  ,.p_bsg_link_in11_tkn_i(GW_IC_LINK_TKN  [11])
  ,.p_bsg_link_in11_d0_o (GW_IC_LINK_D0   [11])
  ,.p_bsg_link_in11_d1_o (GW_IC_LINK_D1   [11])
  ,.p_bsg_link_in11_d2_o (GW_IC_LINK_D2   [11])
  ,.p_bsg_link_in11_d3_o (GW_IC_LINK_D3   [11])
  ,.p_bsg_link_in11_d4_o (GW_IC_LINK_D4   [11])
  ,.p_bsg_link_in11_d5_o (GW_IC_LINK_D5   [11])
  ,.p_bsg_link_in11_d6_o (GW_IC_LINK_D6   [11])
  ,.p_bsg_link_in11_d7_o (GW_IC_LINK_D7   [11])
  ,.p_bsg_link_in11_d8_o (GW_IC_LINK_D8   [11])
                           
  ,.p_bsg_link_in12_clk_o(GW_IC_LINK_CLK  [12])
  ,.p_bsg_link_in12_v_o  (GW_IC_LINK_V    [12])
  ,.p_bsg_link_in12_tkn_i(GW_IC_LINK_TKN  [12])
  ,.p_bsg_link_in12_d0_o (GW_IC_LINK_D0   [12])
  ,.p_bsg_link_in12_d1_o (GW_IC_LINK_D1   [12])
  ,.p_bsg_link_in12_d2_o (GW_IC_LINK_D2   [12])
  ,.p_bsg_link_in12_d3_o (GW_IC_LINK_D3   [12])
  ,.p_bsg_link_in12_d4_o (GW_IC_LINK_D4   [12])
  ,.p_bsg_link_in12_d5_o (GW_IC_LINK_D5   [12])
  ,.p_bsg_link_in12_d6_o (GW_IC_LINK_D6   [12])
  ,.p_bsg_link_in12_d7_o (GW_IC_LINK_D7   [12])
  ,.p_bsg_link_in12_d8_o (GW_IC_LINK_D8   [12])
                           
  ,.p_bsg_link_in13_clk_o(GW_IC_LINK_CLK  [13])
  ,.p_bsg_link_in13_v_o  (GW_IC_LINK_V    [13])
  ,.p_bsg_link_in13_tkn_i(GW_IC_LINK_TKN  [13])
  ,.p_bsg_link_in13_d0_o (GW_IC_LINK_D0   [13])
  ,.p_bsg_link_in13_d1_o (GW_IC_LINK_D1   [13])
  ,.p_bsg_link_in13_d2_o (GW_IC_LINK_D2   [13])
  ,.p_bsg_link_in13_d3_o (GW_IC_LINK_D3   [13])
  ,.p_bsg_link_in13_d4_o (GW_IC_LINK_D4   [13])
  ,.p_bsg_link_in13_d5_o (GW_IC_LINK_D5   [13])
  ,.p_bsg_link_in13_d6_o (GW_IC_LINK_D6   [13])
  ,.p_bsg_link_in13_d7_o (GW_IC_LINK_D7   [13])
  ,.p_bsg_link_in13_d8_o (GW_IC_LINK_D8   [13])
                           
  ,.p_bsg_link_in14_clk_o(GW_IC_LINK_CLK  [14])
  ,.p_bsg_link_in14_v_o  (GW_IC_LINK_V    [14])
  ,.p_bsg_link_in14_tkn_i(GW_IC_LINK_TKN  [14])
  ,.p_bsg_link_in14_d0_o (GW_IC_LINK_D0   [14])
  ,.p_bsg_link_in14_d1_o (GW_IC_LINK_D1   [14])
  ,.p_bsg_link_in14_d2_o (GW_IC_LINK_D2   [14])
  ,.p_bsg_link_in14_d3_o (GW_IC_LINK_D3   [14])
  ,.p_bsg_link_in14_d4_o (GW_IC_LINK_D4   [14])
  ,.p_bsg_link_in14_d5_o (GW_IC_LINK_D5   [14])
  ,.p_bsg_link_in14_d6_o (GW_IC_LINK_D6   [14])
  ,.p_bsg_link_in14_d7_o (GW_IC_LINK_D7   [14])
  ,.p_bsg_link_in14_d8_o (GW_IC_LINK_D8   [14])
                          
  ,.p_bsg_link_in15_clk_o(GW_IC_LINK_CLK  [15])
  ,.p_bsg_link_in15_v_o  (GW_IC_LINK_V    [15])
  ,.p_bsg_link_in15_tkn_i(GW_IC_LINK_TKN  [15])
  ,.p_bsg_link_in15_d0_o (GW_IC_LINK_D0   [15])
  ,.p_bsg_link_in15_d1_o (GW_IC_LINK_D1   [15])
  ,.p_bsg_link_in15_d2_o (GW_IC_LINK_D2   [15])
  ,.p_bsg_link_in15_d3_o (GW_IC_LINK_D3   [15])
  ,.p_bsg_link_in15_d4_o (GW_IC_LINK_D4   [15])
  ,.p_bsg_link_in15_d5_o (GW_IC_LINK_D5   [15])
  ,.p_bsg_link_in15_d6_o (GW_IC_LINK_D6   [15])
  ,.p_bsg_link_in15_d7_o (GW_IC_LINK_D7   [15])
  ,.p_bsg_link_in15_d8_o (GW_IC_LINK_D8   [15])
                           
  ,.p_bsg_link_in16_clk_o(GW_IC_LINK_CLK  [16])
  ,.p_bsg_link_in16_v_o  (GW_IC_LINK_V    [16])
  ,.p_bsg_link_in16_tkn_i(GW_IC_LINK_TKN  [16])
  ,.p_bsg_link_in16_d0_o (GW_IC_LINK_D0   [16])
  ,.p_bsg_link_in16_d1_o (GW_IC_LINK_D1   [16])
  ,.p_bsg_link_in16_d2_o (GW_IC_LINK_D2   [16])
  ,.p_bsg_link_in16_d3_o (GW_IC_LINK_D3   [16])
  ,.p_bsg_link_in16_d4_o (GW_IC_LINK_D4   [16])
  ,.p_bsg_link_in16_d5_o (GW_IC_LINK_D5   [16])
  ,.p_bsg_link_in16_d6_o (GW_IC_LINK_D6   [16])
  ,.p_bsg_link_in16_d7_o (GW_IC_LINK_D7   [16])
  ,.p_bsg_link_in16_d8_o (GW_IC_LINK_D8   [16])
                           
  ,.p_bsg_link_in17_clk_o(GW_IC_LINK_CLK  [17])
  ,.p_bsg_link_in17_v_o  (GW_IC_LINK_V    [17])
  ,.p_bsg_link_in17_tkn_i(GW_IC_LINK_TKN  [17])
  ,.p_bsg_link_in17_d0_o (GW_IC_LINK_D0   [17])
  ,.p_bsg_link_in17_d1_o (GW_IC_LINK_D1   [17])
  ,.p_bsg_link_in17_d2_o (GW_IC_LINK_D2   [17])
  ,.p_bsg_link_in17_d3_o (GW_IC_LINK_D3   [17])
  ,.p_bsg_link_in17_d4_o (GW_IC_LINK_D4   [17])
  ,.p_bsg_link_in17_d5_o (GW_IC_LINK_D5   [17])
  ,.p_bsg_link_in17_d6_o (GW_IC_LINK_D6   [17])
  ,.p_bsg_link_in17_d7_o (GW_IC_LINK_D7   [17])
  ,.p_bsg_link_in17_d8_o (GW_IC_LINK_D8   [17])
                           
  ,.p_bsg_link_in18_clk_o(GW_IC_LINK_CLK  [18])
  ,.p_bsg_link_in18_v_o  (GW_IC_LINK_V    [18])
  ,.p_bsg_link_in18_tkn_i(GW_IC_LINK_TKN  [18])
  ,.p_bsg_link_in18_d0_o (GW_IC_LINK_D0   [18])
  ,.p_bsg_link_in18_d1_o (GW_IC_LINK_D1   [18])
  ,.p_bsg_link_in18_d2_o (GW_IC_LINK_D2   [18])
  ,.p_bsg_link_in18_d3_o (GW_IC_LINK_D3   [18])
  ,.p_bsg_link_in18_d4_o (GW_IC_LINK_D4   [18])
  ,.p_bsg_link_in18_d5_o (GW_IC_LINK_D5   [18])
  ,.p_bsg_link_in18_d6_o (GW_IC_LINK_D6   [18])
  ,.p_bsg_link_in18_d7_o (GW_IC_LINK_D7   [18])
  ,.p_bsg_link_in18_d8_o (GW_IC_LINK_D8   [18])
                           
  ,.p_bsg_link_in19_clk_o(GW_IC_LINK_CLK  [19])
  ,.p_bsg_link_in19_v_o  (GW_IC_LINK_V    [19])
  ,.p_bsg_link_in19_tkn_i(GW_IC_LINK_TKN  [19])
  ,.p_bsg_link_in19_d0_o (GW_IC_LINK_D0   [19])
  ,.p_bsg_link_in19_d1_o (GW_IC_LINK_D1   [19])
  ,.p_bsg_link_in19_d2_o (GW_IC_LINK_D2   [19])
  ,.p_bsg_link_in19_d3_o (GW_IC_LINK_D3   [19])
  ,.p_bsg_link_in19_d4_o (GW_IC_LINK_D4   [19])
  ,.p_bsg_link_in19_d5_o (GW_IC_LINK_D5   [19])
  ,.p_bsg_link_in19_d6_o (GW_IC_LINK_D6   [19])
  ,.p_bsg_link_in19_d7_o (GW_IC_LINK_D7   [19])
  ,.p_bsg_link_in19_d8_o (GW_IC_LINK_D8   [19])
  
  ,.p_bsg_link_out0_clk_i  (IC_GW_LINK_CLK  [0])
  ,.p_bsg_link_out0_v_i    (IC_GW_LINK_V    [0])
  ,.p_bsg_link_out0_tkn_o  (IC_GW_LINK_TKN  [0])
  ,.p_bsg_link_out0_d0_i   (IC_GW_LINK_D0   [0])
  ,.p_bsg_link_out0_d1_i   (IC_GW_LINK_D1   [0])
  ,.p_bsg_link_out0_d2_i   (IC_GW_LINK_D2   [0])
  ,.p_bsg_link_out0_d3_i   (IC_GW_LINK_D3   [0])
  ,.p_bsg_link_out0_d4_i   (IC_GW_LINK_D4   [0])
  ,.p_bsg_link_out0_d5_i   (IC_GW_LINK_D5   [0])
  ,.p_bsg_link_out0_d6_i   (IC_GW_LINK_D6   [0])
  ,.p_bsg_link_out0_d7_i   (IC_GW_LINK_D7   [0])
  ,.p_bsg_link_out0_d8_i   (IC_GW_LINK_D8   [0])
                          
  ,.p_bsg_link_out1_clk_i  (IC_GW_LINK_CLK  [1])
  ,.p_bsg_link_out1_v_i    (IC_GW_LINK_V    [1])
  ,.p_bsg_link_out1_tkn_o  (IC_GW_LINK_TKN  [1])
  ,.p_bsg_link_out1_d0_i   (IC_GW_LINK_D0   [1])
  ,.p_bsg_link_out1_d1_i   (IC_GW_LINK_D1   [1])
  ,.p_bsg_link_out1_d2_i   (IC_GW_LINK_D2   [1])
  ,.p_bsg_link_out1_d3_i   (IC_GW_LINK_D3   [1])
  ,.p_bsg_link_out1_d4_i   (IC_GW_LINK_D4   [1])
  ,.p_bsg_link_out1_d5_i   (IC_GW_LINK_D5   [1])
  ,.p_bsg_link_out1_d6_i   (IC_GW_LINK_D6   [1])
  ,.p_bsg_link_out1_d7_i   (IC_GW_LINK_D7   [1])
  ,.p_bsg_link_out1_d8_i   (IC_GW_LINK_D8   [1])
                          
  ,.p_bsg_link_out2_clk_i  (IC_GW_LINK_CLK  [2])
  ,.p_bsg_link_out2_v_i    (IC_GW_LINK_V    [2])
  ,.p_bsg_link_out2_tkn_o  (IC_GW_LINK_TKN  [2])
  ,.p_bsg_link_out2_d0_i   (IC_GW_LINK_D0   [2])
  ,.p_bsg_link_out2_d1_i   (IC_GW_LINK_D1   [2])
  ,.p_bsg_link_out2_d2_i   (IC_GW_LINK_D2   [2])
  ,.p_bsg_link_out2_d3_i   (IC_GW_LINK_D3   [2])
  ,.p_bsg_link_out2_d4_i   (IC_GW_LINK_D4   [2])
  ,.p_bsg_link_out2_d5_i   (IC_GW_LINK_D5   [2])
  ,.p_bsg_link_out2_d6_i   (IC_GW_LINK_D6   [2])
  ,.p_bsg_link_out2_d7_i   (IC_GW_LINK_D7   [2])
  ,.p_bsg_link_out2_d8_i   (IC_GW_LINK_D8   [2])
                          
  ,.p_bsg_link_out3_clk_i  (IC_GW_LINK_CLK  [3])
  ,.p_bsg_link_out3_v_i    (IC_GW_LINK_V    [3])
  ,.p_bsg_link_out3_tkn_o  (IC_GW_LINK_TKN  [3])
  ,.p_bsg_link_out3_d0_i   (IC_GW_LINK_D0   [3])
  ,.p_bsg_link_out3_d1_i   (IC_GW_LINK_D1   [3])
  ,.p_bsg_link_out3_d2_i   (IC_GW_LINK_D2   [3])
  ,.p_bsg_link_out3_d3_i   (IC_GW_LINK_D3   [3])
  ,.p_bsg_link_out3_d4_i   (IC_GW_LINK_D4   [3])
  ,.p_bsg_link_out3_d5_i   (IC_GW_LINK_D5   [3])
  ,.p_bsg_link_out3_d6_i   (IC_GW_LINK_D6   [3])
  ,.p_bsg_link_out3_d7_i   (IC_GW_LINK_D7   [3])
  ,.p_bsg_link_out3_d8_i   (IC_GW_LINK_D8   [3])
                          
  ,.p_bsg_link_out4_clk_i  (IC_GW_LINK_CLK  [4])
  ,.p_bsg_link_out4_v_i    (IC_GW_LINK_V    [4])
  ,.p_bsg_link_out4_tkn_o  (IC_GW_LINK_TKN  [4])
  ,.p_bsg_link_out4_d0_i   (IC_GW_LINK_D0   [4])
  ,.p_bsg_link_out4_d1_i   (IC_GW_LINK_D1   [4])
  ,.p_bsg_link_out4_d2_i   (IC_GW_LINK_D2   [4])
  ,.p_bsg_link_out4_d3_i   (IC_GW_LINK_D3   [4])
  ,.p_bsg_link_out4_d4_i   (IC_GW_LINK_D4   [4])
  ,.p_bsg_link_out4_d5_i   (IC_GW_LINK_D5   [4])
  ,.p_bsg_link_out4_d6_i   (IC_GW_LINK_D6   [4])
  ,.p_bsg_link_out4_d7_i   (IC_GW_LINK_D7   [4])
  ,.p_bsg_link_out4_d8_i   (IC_GW_LINK_D8   [4])
                          
  ,.p_bsg_link_out5_clk_i  (IC_GW_LINK_CLK  [5])
  ,.p_bsg_link_out5_v_i    (IC_GW_LINK_V    [5])
  ,.p_bsg_link_out5_tkn_o  (IC_GW_LINK_TKN  [5])
  ,.p_bsg_link_out5_d0_i   (IC_GW_LINK_D0   [5])
  ,.p_bsg_link_out5_d1_i   (IC_GW_LINK_D1   [5])
  ,.p_bsg_link_out5_d2_i   (IC_GW_LINK_D2   [5])
  ,.p_bsg_link_out5_d3_i   (IC_GW_LINK_D3   [5])
  ,.p_bsg_link_out5_d4_i   (IC_GW_LINK_D4   [5])
  ,.p_bsg_link_out5_d5_i   (IC_GW_LINK_D5   [5])
  ,.p_bsg_link_out5_d6_i   (IC_GW_LINK_D6   [5])
  ,.p_bsg_link_out5_d7_i   (IC_GW_LINK_D7   [5])
  ,.p_bsg_link_out5_d8_i   (IC_GW_LINK_D8   [5])
                           
  ,.p_bsg_link_out6_clk_i  (IC_GW_LINK_CLK  [6])
  ,.p_bsg_link_out6_v_i    (IC_GW_LINK_V    [6])
  ,.p_bsg_link_out6_tkn_o  (IC_GW_LINK_TKN  [6])
  ,.p_bsg_link_out6_d0_i   (IC_GW_LINK_D0   [6])
  ,.p_bsg_link_out6_d1_i   (IC_GW_LINK_D1   [6])
  ,.p_bsg_link_out6_d2_i   (IC_GW_LINK_D2   [6])
  ,.p_bsg_link_out6_d3_i   (IC_GW_LINK_D3   [6])
  ,.p_bsg_link_out6_d4_i   (IC_GW_LINK_D4   [6])
  ,.p_bsg_link_out6_d5_i   (IC_GW_LINK_D5   [6])
  ,.p_bsg_link_out6_d6_i   (IC_GW_LINK_D6   [6])
  ,.p_bsg_link_out6_d7_i   (IC_GW_LINK_D7   [6])
  ,.p_bsg_link_out6_d8_i   (IC_GW_LINK_D8   [6])
                           
  ,.p_bsg_link_out7_clk_i  (IC_GW_LINK_CLK  [7])
  ,.p_bsg_link_out7_v_i    (IC_GW_LINK_V    [7])
  ,.p_bsg_link_out7_tkn_o  (IC_GW_LINK_TKN  [7])
  ,.p_bsg_link_out7_d0_i   (IC_GW_LINK_D0   [7])
  ,.p_bsg_link_out7_d1_i   (IC_GW_LINK_D1   [7])
  ,.p_bsg_link_out7_d2_i   (IC_GW_LINK_D2   [7])
  ,.p_bsg_link_out7_d3_i   (IC_GW_LINK_D3   [7])
  ,.p_bsg_link_out7_d4_i   (IC_GW_LINK_D4   [7])
  ,.p_bsg_link_out7_d5_i   (IC_GW_LINK_D5   [7])
  ,.p_bsg_link_out7_d6_i   (IC_GW_LINK_D6   [7])
  ,.p_bsg_link_out7_d7_i   (IC_GW_LINK_D7   [7])
  ,.p_bsg_link_out7_d8_i   (IC_GW_LINK_D8   [7])
                           
  ,.p_bsg_link_out8_clk_i  (IC_GW_LINK_CLK  [8])
  ,.p_bsg_link_out8_v_i    (IC_GW_LINK_V    [8])
  ,.p_bsg_link_out8_tkn_o  (IC_GW_LINK_TKN  [8])
  ,.p_bsg_link_out8_d0_i   (IC_GW_LINK_D0   [8])
  ,.p_bsg_link_out8_d1_i   (IC_GW_LINK_D1   [8])
  ,.p_bsg_link_out8_d2_i   (IC_GW_LINK_D2   [8])
  ,.p_bsg_link_out8_d3_i   (IC_GW_LINK_D3   [8])
  ,.p_bsg_link_out8_d4_i   (IC_GW_LINK_D4   [8])
  ,.p_bsg_link_out8_d5_i   (IC_GW_LINK_D5   [8])
  ,.p_bsg_link_out8_d6_i   (IC_GW_LINK_D6   [8])
  ,.p_bsg_link_out8_d7_i   (IC_GW_LINK_D7   [8])
  ,.p_bsg_link_out8_d8_i   (IC_GW_LINK_D8   [8])
                           
  ,.p_bsg_link_out9_clk_i  (IC_GW_LINK_CLK  [9])
  ,.p_bsg_link_out9_v_i    (IC_GW_LINK_V    [9])
  ,.p_bsg_link_out9_tkn_o  (IC_GW_LINK_TKN  [9])
  ,.p_bsg_link_out9_d0_i   (IC_GW_LINK_D0   [9])
  ,.p_bsg_link_out9_d1_i   (IC_GW_LINK_D1   [9])
  ,.p_bsg_link_out9_d2_i   (IC_GW_LINK_D2   [9])
  ,.p_bsg_link_out9_d3_i   (IC_GW_LINK_D3   [9])
  ,.p_bsg_link_out9_d4_i   (IC_GW_LINK_D4   [9])
  ,.p_bsg_link_out9_d5_i   (IC_GW_LINK_D5   [9])
  ,.p_bsg_link_out9_d6_i   (IC_GW_LINK_D6   [9])
  ,.p_bsg_link_out9_d7_i   (IC_GW_LINK_D7   [9])
  ,.p_bsg_link_out9_d8_i   (IC_GW_LINK_D8   [9])
                          
  ,.p_bsg_link_out10_clk_i (IC_GW_LINK_CLK  [10])
  ,.p_bsg_link_out10_v_i   (IC_GW_LINK_V    [10])
  ,.p_bsg_link_out10_tkn_o (IC_GW_LINK_TKN  [10])
  ,.p_bsg_link_out10_d0_i  (IC_GW_LINK_D0   [10])
  ,.p_bsg_link_out10_d1_i  (IC_GW_LINK_D1   [10])
  ,.p_bsg_link_out10_d2_i  (IC_GW_LINK_D2   [10])
  ,.p_bsg_link_out10_d3_i  (IC_GW_LINK_D3   [10])
  ,.p_bsg_link_out10_d4_i  (IC_GW_LINK_D4   [10])
  ,.p_bsg_link_out10_d5_i  (IC_GW_LINK_D5   [10])
  ,.p_bsg_link_out10_d6_i  (IC_GW_LINK_D6   [10])
  ,.p_bsg_link_out10_d7_i  (IC_GW_LINK_D7   [10])
  ,.p_bsg_link_out10_d8_i  (IC_GW_LINK_D8   [10])
                           
  ,.p_bsg_link_out11_clk_i (IC_GW_LINK_CLK  [11])
  ,.p_bsg_link_out11_v_i   (IC_GW_LINK_V    [11])
  ,.p_bsg_link_out11_tkn_o (IC_GW_LINK_TKN  [11])
  ,.p_bsg_link_out11_d0_i  (IC_GW_LINK_D0   [11])
  ,.p_bsg_link_out11_d1_i  (IC_GW_LINK_D1   [11])
  ,.p_bsg_link_out11_d2_i  (IC_GW_LINK_D2   [11])
  ,.p_bsg_link_out11_d3_i  (IC_GW_LINK_D3   [11])
  ,.p_bsg_link_out11_d4_i  (IC_GW_LINK_D4   [11])
  ,.p_bsg_link_out11_d5_i  (IC_GW_LINK_D5   [11])
  ,.p_bsg_link_out11_d6_i  (IC_GW_LINK_D6   [11])
  ,.p_bsg_link_out11_d7_i  (IC_GW_LINK_D7   [11])
  ,.p_bsg_link_out11_d8_i  (IC_GW_LINK_D8   [11])
                           
  ,.p_bsg_link_out12_clk_i (IC_GW_LINK_CLK  [12])
  ,.p_bsg_link_out12_v_i   (IC_GW_LINK_V    [12])
  ,.p_bsg_link_out12_tkn_o (IC_GW_LINK_TKN  [12])
  ,.p_bsg_link_out12_d0_i  (IC_GW_LINK_D0   [12])
  ,.p_bsg_link_out12_d1_i  (IC_GW_LINK_D1   [12])
  ,.p_bsg_link_out12_d2_i  (IC_GW_LINK_D2   [12])
  ,.p_bsg_link_out12_d3_i  (IC_GW_LINK_D3   [12])
  ,.p_bsg_link_out12_d4_i  (IC_GW_LINK_D4   [12])
  ,.p_bsg_link_out12_d5_i  (IC_GW_LINK_D5   [12])
  ,.p_bsg_link_out12_d6_i  (IC_GW_LINK_D6   [12])
  ,.p_bsg_link_out12_d7_i  (IC_GW_LINK_D7   [12])
  ,.p_bsg_link_out12_d8_i  (IC_GW_LINK_D8   [12])
                           
  ,.p_bsg_link_out13_clk_i (IC_GW_LINK_CLK  [13])
  ,.p_bsg_link_out13_v_i   (IC_GW_LINK_V    [13])
  ,.p_bsg_link_out13_tkn_o (IC_GW_LINK_TKN  [13])
  ,.p_bsg_link_out13_d0_i  (IC_GW_LINK_D0   [13])
  ,.p_bsg_link_out13_d1_i  (IC_GW_LINK_D1   [13])
  ,.p_bsg_link_out13_d2_i  (IC_GW_LINK_D2   [13])
  ,.p_bsg_link_out13_d3_i  (IC_GW_LINK_D3   [13])
  ,.p_bsg_link_out13_d4_i  (IC_GW_LINK_D4   [13])
  ,.p_bsg_link_out13_d5_i  (IC_GW_LINK_D5   [13])
  ,.p_bsg_link_out13_d6_i  (IC_GW_LINK_D6   [13])
  ,.p_bsg_link_out13_d7_i  (IC_GW_LINK_D7   [13])
  ,.p_bsg_link_out13_d8_i  (IC_GW_LINK_D8   [13])
                           
  ,.p_bsg_link_out14_clk_i (IC_GW_LINK_CLK  [14])
  ,.p_bsg_link_out14_v_i   (IC_GW_LINK_V    [14])
  ,.p_bsg_link_out14_tkn_o (IC_GW_LINK_TKN  [14])
  ,.p_bsg_link_out14_d0_i  (IC_GW_LINK_D0   [14])
  ,.p_bsg_link_out14_d1_i  (IC_GW_LINK_D1   [14])
  ,.p_bsg_link_out14_d2_i  (IC_GW_LINK_D2   [14])
  ,.p_bsg_link_out14_d3_i  (IC_GW_LINK_D3   [14])
  ,.p_bsg_link_out14_d4_i  (IC_GW_LINK_D4   [14])
  ,.p_bsg_link_out14_d5_i  (IC_GW_LINK_D5   [14])
  ,.p_bsg_link_out14_d6_i  (IC_GW_LINK_D6   [14])
  ,.p_bsg_link_out14_d7_i  (IC_GW_LINK_D7   [14])
  ,.p_bsg_link_out14_d8_i  (IC_GW_LINK_D8   [14])
                          
  ,.p_bsg_link_out15_clk_i (IC_GW_LINK_CLK  [15])
  ,.p_bsg_link_out15_v_i   (IC_GW_LINK_V    [15])
  ,.p_bsg_link_out15_tkn_o (IC_GW_LINK_TKN  [15])
  ,.p_bsg_link_out15_d0_i  (IC_GW_LINK_D0   [15])
  ,.p_bsg_link_out15_d1_i  (IC_GW_LINK_D1   [15])
  ,.p_bsg_link_out15_d2_i  (IC_GW_LINK_D2   [15])
  ,.p_bsg_link_out15_d3_i  (IC_GW_LINK_D3   [15])
  ,.p_bsg_link_out15_d4_i  (IC_GW_LINK_D4   [15])
  ,.p_bsg_link_out15_d5_i  (IC_GW_LINK_D5   [15])
  ,.p_bsg_link_out15_d6_i  (IC_GW_LINK_D6   [15])
  ,.p_bsg_link_out15_d7_i  (IC_GW_LINK_D7   [15])
  ,.p_bsg_link_out15_d8_i  (IC_GW_LINK_D8   [15])
                           
  ,.p_bsg_link_out16_clk_i (IC_GW_LINK_CLK  [16])
  ,.p_bsg_link_out16_v_i   (IC_GW_LINK_V    [16])
  ,.p_bsg_link_out16_tkn_o (IC_GW_LINK_TKN  [16])
  ,.p_bsg_link_out16_d0_i  (IC_GW_LINK_D0   [16])
  ,.p_bsg_link_out16_d1_i  (IC_GW_LINK_D1   [16])
  ,.p_bsg_link_out16_d2_i  (IC_GW_LINK_D2   [16])
  ,.p_bsg_link_out16_d3_i  (IC_GW_LINK_D3   [16])
  ,.p_bsg_link_out16_d4_i  (IC_GW_LINK_D4   [16])
  ,.p_bsg_link_out16_d5_i  (IC_GW_LINK_D5   [16])
  ,.p_bsg_link_out16_d6_i  (IC_GW_LINK_D6   [16])
  ,.p_bsg_link_out16_d7_i  (IC_GW_LINK_D7   [16])
  ,.p_bsg_link_out16_d8_i  (IC_GW_LINK_D8   [16])
                           
  ,.p_bsg_link_out17_clk_i (IC_GW_LINK_CLK  [17])
  ,.p_bsg_link_out17_v_i   (IC_GW_LINK_V    [17])
  ,.p_bsg_link_out17_tkn_o (IC_GW_LINK_TKN  [17])
  ,.p_bsg_link_out17_d0_i  (IC_GW_LINK_D0   [17])
  ,.p_bsg_link_out17_d1_i  (IC_GW_LINK_D1   [17])
  ,.p_bsg_link_out17_d2_i  (IC_GW_LINK_D2   [17])
  ,.p_bsg_link_out17_d3_i  (IC_GW_LINK_D3   [17])
  ,.p_bsg_link_out17_d4_i  (IC_GW_LINK_D4   [17])
  ,.p_bsg_link_out17_d5_i  (IC_GW_LINK_D5   [17])
  ,.p_bsg_link_out17_d6_i  (IC_GW_LINK_D6   [17])
  ,.p_bsg_link_out17_d7_i  (IC_GW_LINK_D7   [17])
  ,.p_bsg_link_out17_d8_i  (IC_GW_LINK_D8   [17])
                           
  ,.p_bsg_link_out18_clk_i (IC_GW_LINK_CLK  [18])
  ,.p_bsg_link_out18_v_i   (IC_GW_LINK_V    [18])
  ,.p_bsg_link_out18_tkn_o (IC_GW_LINK_TKN  [18])
  ,.p_bsg_link_out18_d0_i  (IC_GW_LINK_D0   [18])
  ,.p_bsg_link_out18_d1_i  (IC_GW_LINK_D1   [18])
  ,.p_bsg_link_out18_d2_i  (IC_GW_LINK_D2   [18])
  ,.p_bsg_link_out18_d3_i  (IC_GW_LINK_D3   [18])
  ,.p_bsg_link_out18_d4_i  (IC_GW_LINK_D4   [18])
  ,.p_bsg_link_out18_d5_i  (IC_GW_LINK_D5   [18])
  ,.p_bsg_link_out18_d6_i  (IC_GW_LINK_D6   [18])
  ,.p_bsg_link_out18_d7_i  (IC_GW_LINK_D7   [18])
  ,.p_bsg_link_out18_d8_i  (IC_GW_LINK_D8   [18])
                           
  ,.p_bsg_link_out19_clk_i (IC_GW_LINK_CLK  [19])
  ,.p_bsg_link_out19_v_i   (IC_GW_LINK_V    [19])
  ,.p_bsg_link_out19_tkn_o (IC_GW_LINK_TKN  [19])
  ,.p_bsg_link_out19_d0_i  (IC_GW_LINK_D0   [19])
  ,.p_bsg_link_out19_d1_i  (IC_GW_LINK_D1   [19])
  ,.p_bsg_link_out19_d2_i  (IC_GW_LINK_D2   [19])
  ,.p_bsg_link_out19_d3_i  (IC_GW_LINK_D3   [19])
  ,.p_bsg_link_out19_d4_i  (IC_GW_LINK_D4   [19])
  ,.p_bsg_link_out19_d5_i  (IC_GW_LINK_D5   [19])
  ,.p_bsg_link_out19_d6_i  (IC_GW_LINK_D6   [19])
  ,.p_bsg_link_out19_d7_i  (IC_GW_LINK_D7   [19])
  ,.p_bsg_link_out19_d8_i  (IC_GW_LINK_D8   [19])

  ,.p_bsg_tag_clk_o       (GW_TAG_CLKO)
  ,.p_bsg_tag_en_o        (GW_TAG_EN)
  ,.p_bsg_tag_data_o      (GW_TAG_DATAO)
  ,.p_bsg_tag_clk_i       ()
  ,.p_bsg_tag_data_i      ()

  ,.p_clk_A_o             (GW_CLKA)
  ,.p_clk_B_o             (GW_CLKB)
  ,.p_clk_C_o             (GW_CLKC)

  ,.p_clk_i               (IC_CLKO)

  ,.p_sel_0_o             (GW_SEL0)
  ,.p_sel_1_o             (GW_SEL1)
  ,.p_sel_2_o             (GW_SEL2)

  ,.p_clk_async_reset_o   (GW_CLK_RESET)
  ,.p_core_async_reset_o  (GW_CORE_RESET)

  ,.p_misc_i              ()
  );

  //
  // ASIC SOCKET
  //

  bsg_chip IC
  (.p_bsg_link_in0_clk_i  (GW_IC_LINK_CLK  [0])
  ,.p_bsg_link_in0_v_i    (GW_IC_LINK_V    [0])
  ,.p_bsg_link_in0_tkn_o  (GW_IC_LINK_TKN  [0])
  ,.p_bsg_link_in0_d0_i   (GW_IC_LINK_D0   [0])
  ,.p_bsg_link_in0_d1_i   (GW_IC_LINK_D1   [0])
  ,.p_bsg_link_in0_d2_i   (GW_IC_LINK_D2   [0])
  ,.p_bsg_link_in0_d3_i   (GW_IC_LINK_D3   [0])
  ,.p_bsg_link_in0_d4_i   (GW_IC_LINK_D4   [0])
  ,.p_bsg_link_in0_d5_i   (GW_IC_LINK_D5   [0])
  ,.p_bsg_link_in0_d6_i   (GW_IC_LINK_D6   [0])
  ,.p_bsg_link_in0_d7_i   (GW_IC_LINK_D7   [0])
  ,.p_bsg_link_in0_d8_i   (GW_IC_LINK_D8   [0])
                          
  ,.p_bsg_link_in1_clk_i  (GW_IC_LINK_CLK  [1])
  ,.p_bsg_link_in1_v_i    (GW_IC_LINK_V    [1])
  ,.p_bsg_link_in1_tkn_o  (GW_IC_LINK_TKN  [1])
  ,.p_bsg_link_in1_d0_i   (GW_IC_LINK_D0   [1])
  ,.p_bsg_link_in1_d1_i   (GW_IC_LINK_D1   [1])
  ,.p_bsg_link_in1_d2_i   (GW_IC_LINK_D2   [1])
  ,.p_bsg_link_in1_d3_i   (GW_IC_LINK_D3   [1])
  ,.p_bsg_link_in1_d4_i   (GW_IC_LINK_D4   [1])
  ,.p_bsg_link_in1_d5_i   (GW_IC_LINK_D5   [1])
  ,.p_bsg_link_in1_d6_i   (GW_IC_LINK_D6   [1])
  ,.p_bsg_link_in1_d7_i   (GW_IC_LINK_D7   [1])
  ,.p_bsg_link_in1_d8_i   (GW_IC_LINK_D8   [1])
                          
  ,.p_bsg_link_in2_clk_i  (GW_IC_LINK_CLK  [2])
  ,.p_bsg_link_in2_v_i    (GW_IC_LINK_V    [2])
  ,.p_bsg_link_in2_tkn_o  (GW_IC_LINK_TKN  [2])
  ,.p_bsg_link_in2_d0_i   (GW_IC_LINK_D0   [2])
  ,.p_bsg_link_in2_d1_i   (GW_IC_LINK_D1   [2])
  ,.p_bsg_link_in2_d2_i   (GW_IC_LINK_D2   [2])
  ,.p_bsg_link_in2_d3_i   (GW_IC_LINK_D3   [2])
  ,.p_bsg_link_in2_d4_i   (GW_IC_LINK_D4   [2])
  ,.p_bsg_link_in2_d5_i   (GW_IC_LINK_D5   [2])
  ,.p_bsg_link_in2_d6_i   (GW_IC_LINK_D6   [2])
  ,.p_bsg_link_in2_d7_i   (GW_IC_LINK_D7   [2])
  ,.p_bsg_link_in2_d8_i   (GW_IC_LINK_D8   [2])
                          
  ,.p_bsg_link_in3_clk_i  (GW_IC_LINK_CLK  [3])
  ,.p_bsg_link_in3_v_i    (GW_IC_LINK_V    [3])
  ,.p_bsg_link_in3_tkn_o  (GW_IC_LINK_TKN  [3])
  ,.p_bsg_link_in3_d0_i   (GW_IC_LINK_D0   [3])
  ,.p_bsg_link_in3_d1_i   (GW_IC_LINK_D1   [3])
  ,.p_bsg_link_in3_d2_i   (GW_IC_LINK_D2   [3])
  ,.p_bsg_link_in3_d3_i   (GW_IC_LINK_D3   [3])
  ,.p_bsg_link_in3_d4_i   (GW_IC_LINK_D4   [3])
  ,.p_bsg_link_in3_d5_i   (GW_IC_LINK_D5   [3])
  ,.p_bsg_link_in3_d6_i   (GW_IC_LINK_D6   [3])
  ,.p_bsg_link_in3_d7_i   (GW_IC_LINK_D7   [3])
  ,.p_bsg_link_in3_d8_i   (GW_IC_LINK_D8   [3])
                          
  ,.p_bsg_link_in4_clk_i  (GW_IC_LINK_CLK  [4])
  ,.p_bsg_link_in4_v_i    (GW_IC_LINK_V    [4])
  ,.p_bsg_link_in4_tkn_o  (GW_IC_LINK_TKN  [4])
  ,.p_bsg_link_in4_d0_i   (GW_IC_LINK_D0   [4])
  ,.p_bsg_link_in4_d1_i   (GW_IC_LINK_D1   [4])
  ,.p_bsg_link_in4_d2_i   (GW_IC_LINK_D2   [4])
  ,.p_bsg_link_in4_d3_i   (GW_IC_LINK_D3   [4])
  ,.p_bsg_link_in4_d4_i   (GW_IC_LINK_D4   [4])
  ,.p_bsg_link_in4_d5_i   (GW_IC_LINK_D5   [4])
  ,.p_bsg_link_in4_d6_i   (GW_IC_LINK_D6   [4])
  ,.p_bsg_link_in4_d7_i   (GW_IC_LINK_D7   [4])
  ,.p_bsg_link_in4_d8_i   (GW_IC_LINK_D8   [4])
                          
  ,.p_bsg_link_in5_clk_i  (GW_IC_LINK_CLK  [5])
  ,.p_bsg_link_in5_v_i    (GW_IC_LINK_V    [5])
  ,.p_bsg_link_in5_tkn_o  (GW_IC_LINK_TKN  [5])
  ,.p_bsg_link_in5_d0_i   (GW_IC_LINK_D0   [5])
  ,.p_bsg_link_in5_d1_i   (GW_IC_LINK_D1   [5])
  ,.p_bsg_link_in5_d2_i   (GW_IC_LINK_D2   [5])
  ,.p_bsg_link_in5_d3_i   (GW_IC_LINK_D3   [5])
  ,.p_bsg_link_in5_d4_i   (GW_IC_LINK_D4   [5])
  ,.p_bsg_link_in5_d5_i   (GW_IC_LINK_D5   [5])
  ,.p_bsg_link_in5_d6_i   (GW_IC_LINK_D6   [5])
  ,.p_bsg_link_in5_d7_i   (GW_IC_LINK_D7   [5])
  ,.p_bsg_link_in5_d8_i   (GW_IC_LINK_D8   [5])
                           
  ,.p_bsg_link_in6_clk_i  (GW_IC_LINK_CLK  [6])
  ,.p_bsg_link_in6_v_i    (GW_IC_LINK_V    [6])
  ,.p_bsg_link_in6_tkn_o  (GW_IC_LINK_TKN  [6])
  ,.p_bsg_link_in6_d0_i   (GW_IC_LINK_D0   [6])
  ,.p_bsg_link_in6_d1_i   (GW_IC_LINK_D1   [6])
  ,.p_bsg_link_in6_d2_i   (GW_IC_LINK_D2   [6])
  ,.p_bsg_link_in6_d3_i   (GW_IC_LINK_D3   [6])
  ,.p_bsg_link_in6_d4_i   (GW_IC_LINK_D4   [6])
  ,.p_bsg_link_in6_d5_i   (GW_IC_LINK_D5   [6])
  ,.p_bsg_link_in6_d6_i   (GW_IC_LINK_D6   [6])
  ,.p_bsg_link_in6_d7_i   (GW_IC_LINK_D7   [6])
  ,.p_bsg_link_in6_d8_i   (GW_IC_LINK_D8   [6])
                           
  ,.p_bsg_link_in7_clk_i  (GW_IC_LINK_CLK  [7])
  ,.p_bsg_link_in7_v_i    (GW_IC_LINK_V    [7])
  ,.p_bsg_link_in7_tkn_o  (GW_IC_LINK_TKN  [7])
  ,.p_bsg_link_in7_d0_i   (GW_IC_LINK_D0   [7])
  ,.p_bsg_link_in7_d1_i   (GW_IC_LINK_D1   [7])
  ,.p_bsg_link_in7_d2_i   (GW_IC_LINK_D2   [7])
  ,.p_bsg_link_in7_d3_i   (GW_IC_LINK_D3   [7])
  ,.p_bsg_link_in7_d4_i   (GW_IC_LINK_D4   [7])
  ,.p_bsg_link_in7_d5_i   (GW_IC_LINK_D5   [7])
  ,.p_bsg_link_in7_d6_i   (GW_IC_LINK_D6   [7])
  ,.p_bsg_link_in7_d7_i   (GW_IC_LINK_D7   [7])
  ,.p_bsg_link_in7_d8_i   (GW_IC_LINK_D8   [7])
                           
  ,.p_bsg_link_in8_clk_i  (GW_IC_LINK_CLK  [8])
  ,.p_bsg_link_in8_v_i    (GW_IC_LINK_V    [8])
  ,.p_bsg_link_in8_tkn_o  (GW_IC_LINK_TKN  [8])
  ,.p_bsg_link_in8_d0_i   (GW_IC_LINK_D0   [8])
  ,.p_bsg_link_in8_d1_i   (GW_IC_LINK_D1   [8])
  ,.p_bsg_link_in8_d2_i   (GW_IC_LINK_D2   [8])
  ,.p_bsg_link_in8_d3_i   (GW_IC_LINK_D3   [8])
  ,.p_bsg_link_in8_d4_i   (GW_IC_LINK_D4   [8])
  ,.p_bsg_link_in8_d5_i   (GW_IC_LINK_D5   [8])
  ,.p_bsg_link_in8_d6_i   (GW_IC_LINK_D6   [8])
  ,.p_bsg_link_in8_d7_i   (GW_IC_LINK_D7   [8])
  ,.p_bsg_link_in8_d8_i   (GW_IC_LINK_D8   [8])
                           
  ,.p_bsg_link_in9_clk_i  (GW_IC_LINK_CLK  [9])
  ,.p_bsg_link_in9_v_i    (GW_IC_LINK_V    [9])
  ,.p_bsg_link_in9_tkn_o  (GW_IC_LINK_TKN  [9])
  ,.p_bsg_link_in9_d0_i   (GW_IC_LINK_D0   [9])
  ,.p_bsg_link_in9_d1_i   (GW_IC_LINK_D1   [9])
  ,.p_bsg_link_in9_d2_i   (GW_IC_LINK_D2   [9])
  ,.p_bsg_link_in9_d3_i   (GW_IC_LINK_D3   [9])
  ,.p_bsg_link_in9_d4_i   (GW_IC_LINK_D4   [9])
  ,.p_bsg_link_in9_d5_i   (GW_IC_LINK_D5   [9])
  ,.p_bsg_link_in9_d6_i   (GW_IC_LINK_D6   [9])
  ,.p_bsg_link_in9_d7_i   (GW_IC_LINK_D7   [9])
  ,.p_bsg_link_in9_d8_i   (GW_IC_LINK_D8   [9])
                          
  ,.p_bsg_link_in10_clk_i (GW_IC_LINK_CLK  [10])
  ,.p_bsg_link_in10_v_i   (GW_IC_LINK_V    [10])
  ,.p_bsg_link_in10_tkn_o (GW_IC_LINK_TKN  [10])
  ,.p_bsg_link_in10_d0_i  (GW_IC_LINK_D0   [10])
  ,.p_bsg_link_in10_d1_i  (GW_IC_LINK_D1   [10])
  ,.p_bsg_link_in10_d2_i  (GW_IC_LINK_D2   [10])
  ,.p_bsg_link_in10_d3_i  (GW_IC_LINK_D3   [10])
  ,.p_bsg_link_in10_d4_i  (GW_IC_LINK_D4   [10])
  ,.p_bsg_link_in10_d5_i  (GW_IC_LINK_D5   [10])
  ,.p_bsg_link_in10_d6_i  (GW_IC_LINK_D6   [10])
  ,.p_bsg_link_in10_d7_i  (GW_IC_LINK_D7   [10])
  ,.p_bsg_link_in10_d8_i  (GW_IC_LINK_D8   [10])
                           
  ,.p_bsg_link_in11_clk_i (GW_IC_LINK_CLK  [11])
  ,.p_bsg_link_in11_v_i   (GW_IC_LINK_V    [11])
  ,.p_bsg_link_in11_tkn_o (GW_IC_LINK_TKN  [11])
  ,.p_bsg_link_in11_d0_i  (GW_IC_LINK_D0   [11])
  ,.p_bsg_link_in11_d1_i  (GW_IC_LINK_D1   [11])
  ,.p_bsg_link_in11_d2_i  (GW_IC_LINK_D2   [11])
  ,.p_bsg_link_in11_d3_i  (GW_IC_LINK_D3   [11])
  ,.p_bsg_link_in11_d4_i  (GW_IC_LINK_D4   [11])
  ,.p_bsg_link_in11_d5_i  (GW_IC_LINK_D5   [11])
  ,.p_bsg_link_in11_d6_i  (GW_IC_LINK_D6   [11])
  ,.p_bsg_link_in11_d7_i  (GW_IC_LINK_D7   [11])
  ,.p_bsg_link_in11_d8_i  (GW_IC_LINK_D8   [11])
                           
  ,.p_bsg_link_in12_clk_i (GW_IC_LINK_CLK  [12])
  ,.p_bsg_link_in12_v_i   (GW_IC_LINK_V    [12])
  ,.p_bsg_link_in12_tkn_o (GW_IC_LINK_TKN  [12])
  ,.p_bsg_link_in12_d0_i  (GW_IC_LINK_D0   [12])
  ,.p_bsg_link_in12_d1_i  (GW_IC_LINK_D1   [12])
  ,.p_bsg_link_in12_d2_i  (GW_IC_LINK_D2   [12])
  ,.p_bsg_link_in12_d3_i  (GW_IC_LINK_D3   [12])
  ,.p_bsg_link_in12_d4_i  (GW_IC_LINK_D4   [12])
  ,.p_bsg_link_in12_d5_i  (GW_IC_LINK_D5   [12])
  ,.p_bsg_link_in12_d6_i  (GW_IC_LINK_D6   [12])
  ,.p_bsg_link_in12_d7_i  (GW_IC_LINK_D7   [12])
  ,.p_bsg_link_in12_d8_i  (GW_IC_LINK_D8   [12])
                           
  ,.p_bsg_link_in13_clk_i (GW_IC_LINK_CLK  [13])
  ,.p_bsg_link_in13_v_i   (GW_IC_LINK_V    [13])
  ,.p_bsg_link_in13_tkn_o (GW_IC_LINK_TKN  [13])
  ,.p_bsg_link_in13_d0_i  (GW_IC_LINK_D0   [13])
  ,.p_bsg_link_in13_d1_i  (GW_IC_LINK_D1   [13])
  ,.p_bsg_link_in13_d2_i  (GW_IC_LINK_D2   [13])
  ,.p_bsg_link_in13_d3_i  (GW_IC_LINK_D3   [13])
  ,.p_bsg_link_in13_d4_i  (GW_IC_LINK_D4   [13])
  ,.p_bsg_link_in13_d5_i  (GW_IC_LINK_D5   [13])
  ,.p_bsg_link_in13_d6_i  (GW_IC_LINK_D6   [13])
  ,.p_bsg_link_in13_d7_i  (GW_IC_LINK_D7   [13])
  ,.p_bsg_link_in13_d8_i  (GW_IC_LINK_D8   [13])
                           
  ,.p_bsg_link_in14_clk_i (GW_IC_LINK_CLK  [14])
  ,.p_bsg_link_in14_v_i   (GW_IC_LINK_V    [14])
  ,.p_bsg_link_in14_tkn_o (GW_IC_LINK_TKN  [14])
  ,.p_bsg_link_in14_d0_i  (GW_IC_LINK_D0   [14])
  ,.p_bsg_link_in14_d1_i  (GW_IC_LINK_D1   [14])
  ,.p_bsg_link_in14_d2_i  (GW_IC_LINK_D2   [14])
  ,.p_bsg_link_in14_d3_i  (GW_IC_LINK_D3   [14])
  ,.p_bsg_link_in14_d4_i  (GW_IC_LINK_D4   [14])
  ,.p_bsg_link_in14_d5_i  (GW_IC_LINK_D5   [14])
  ,.p_bsg_link_in14_d6_i  (GW_IC_LINK_D6   [14])
  ,.p_bsg_link_in14_d7_i  (GW_IC_LINK_D7   [14])
  ,.p_bsg_link_in14_d8_i  (GW_IC_LINK_D8   [14])
                          
  ,.p_bsg_link_in15_clk_i (GW_IC_LINK_CLK  [15])
  ,.p_bsg_link_in15_v_i   (GW_IC_LINK_V    [15])
  ,.p_bsg_link_in15_tkn_o (GW_IC_LINK_TKN  [15])
  ,.p_bsg_link_in15_d0_i  (GW_IC_LINK_D0   [15])
  ,.p_bsg_link_in15_d1_i  (GW_IC_LINK_D1   [15])
  ,.p_bsg_link_in15_d2_i  (GW_IC_LINK_D2   [15])
  ,.p_bsg_link_in15_d3_i  (GW_IC_LINK_D3   [15])
  ,.p_bsg_link_in15_d4_i  (GW_IC_LINK_D4   [15])
  ,.p_bsg_link_in15_d5_i  (GW_IC_LINK_D5   [15])
  ,.p_bsg_link_in15_d6_i  (GW_IC_LINK_D6   [15])
  ,.p_bsg_link_in15_d7_i  (GW_IC_LINK_D7   [15])
  ,.p_bsg_link_in15_d8_i  (GW_IC_LINK_D8   [15])
                           
  ,.p_bsg_link_in16_clk_i (GW_IC_LINK_CLK  [16])
  ,.p_bsg_link_in16_v_i   (GW_IC_LINK_V    [16])
  ,.p_bsg_link_in16_tkn_o (GW_IC_LINK_TKN  [16])
  ,.p_bsg_link_in16_d0_i  (GW_IC_LINK_D0   [16])
  ,.p_bsg_link_in16_d1_i  (GW_IC_LINK_D1   [16])
  ,.p_bsg_link_in16_d2_i  (GW_IC_LINK_D2   [16])
  ,.p_bsg_link_in16_d3_i  (GW_IC_LINK_D3   [16])
  ,.p_bsg_link_in16_d4_i  (GW_IC_LINK_D4   [16])
  ,.p_bsg_link_in16_d5_i  (GW_IC_LINK_D5   [16])
  ,.p_bsg_link_in16_d6_i  (GW_IC_LINK_D6   [16])
  ,.p_bsg_link_in16_d7_i  (GW_IC_LINK_D7   [16])
  ,.p_bsg_link_in16_d8_i  (GW_IC_LINK_D8   [16])
                           
  ,.p_bsg_link_in17_clk_i (GW_IC_LINK_CLK  [17])
  ,.p_bsg_link_in17_v_i   (GW_IC_LINK_V    [17])
  ,.p_bsg_link_in17_tkn_o (GW_IC_LINK_TKN  [17])
  ,.p_bsg_link_in17_d0_i  (GW_IC_LINK_D0   [17])
  ,.p_bsg_link_in17_d1_i  (GW_IC_LINK_D1   [17])
  ,.p_bsg_link_in17_d2_i  (GW_IC_LINK_D2   [17])
  ,.p_bsg_link_in17_d3_i  (GW_IC_LINK_D3   [17])
  ,.p_bsg_link_in17_d4_i  (GW_IC_LINK_D4   [17])
  ,.p_bsg_link_in17_d5_i  (GW_IC_LINK_D5   [17])
  ,.p_bsg_link_in17_d6_i  (GW_IC_LINK_D6   [17])
  ,.p_bsg_link_in17_d7_i  (GW_IC_LINK_D7   [17])
  ,.p_bsg_link_in17_d8_i  (GW_IC_LINK_D8   [17])
                           
  ,.p_bsg_link_in18_clk_i (GW_IC_LINK_CLK  [18])
  ,.p_bsg_link_in18_v_i   (GW_IC_LINK_V    [18])
  ,.p_bsg_link_in18_tkn_o (GW_IC_LINK_TKN  [18])
  ,.p_bsg_link_in18_d0_i  (GW_IC_LINK_D0   [18])
  ,.p_bsg_link_in18_d1_i  (GW_IC_LINK_D1   [18])
  ,.p_bsg_link_in18_d2_i  (GW_IC_LINK_D2   [18])
  ,.p_bsg_link_in18_d3_i  (GW_IC_LINK_D3   [18])
  ,.p_bsg_link_in18_d4_i  (GW_IC_LINK_D4   [18])
  ,.p_bsg_link_in18_d5_i  (GW_IC_LINK_D5   [18])
  ,.p_bsg_link_in18_d6_i  (GW_IC_LINK_D6   [18])
  ,.p_bsg_link_in18_d7_i  (GW_IC_LINK_D7   [18])
  ,.p_bsg_link_in18_d8_i  (GW_IC_LINK_D8   [18])
                           
  ,.p_bsg_link_in19_clk_i (GW_IC_LINK_CLK  [19])
  ,.p_bsg_link_in19_v_i   (GW_IC_LINK_V    [19])
  ,.p_bsg_link_in19_tkn_o (GW_IC_LINK_TKN  [19])
  ,.p_bsg_link_in19_d0_i  (GW_IC_LINK_D0   [19])
  ,.p_bsg_link_in19_d1_i  (GW_IC_LINK_D1   [19])
  ,.p_bsg_link_in19_d2_i  (GW_IC_LINK_D2   [19])
  ,.p_bsg_link_in19_d3_i  (GW_IC_LINK_D3   [19])
  ,.p_bsg_link_in19_d4_i  (GW_IC_LINK_D4   [19])
  ,.p_bsg_link_in19_d5_i  (GW_IC_LINK_D5   [19])
  ,.p_bsg_link_in19_d6_i  (GW_IC_LINK_D6   [19])
  ,.p_bsg_link_in19_d7_i  (GW_IC_LINK_D7   [19])
  ,.p_bsg_link_in19_d8_i  (GW_IC_LINK_D8   [19])
                          
  ,.p_bsg_link_out0_clk_o (IC_GW_LINK_CLK  [0])
  ,.p_bsg_link_out0_v_o   (IC_GW_LINK_V    [0])
  ,.p_bsg_link_out0_tkn_i (IC_GW_LINK_TKN  [0])
  ,.p_bsg_link_out0_d0_o  (IC_GW_LINK_D0   [0])
  ,.p_bsg_link_out0_d1_o  (IC_GW_LINK_D1   [0])
  ,.p_bsg_link_out0_d2_o  (IC_GW_LINK_D2   [0])
  ,.p_bsg_link_out0_d3_o  (IC_GW_LINK_D3   [0])
  ,.p_bsg_link_out0_d4_o  (IC_GW_LINK_D4   [0])
  ,.p_bsg_link_out0_d5_o  (IC_GW_LINK_D5   [0])
  ,.p_bsg_link_out0_d6_o  (IC_GW_LINK_D6   [0])
  ,.p_bsg_link_out0_d7_o  (IC_GW_LINK_D7   [0])
  ,.p_bsg_link_out0_d8_o  (IC_GW_LINK_D8   [0])
                          
  ,.p_bsg_link_out1_clk_o (IC_GW_LINK_CLK  [1])
  ,.p_bsg_link_out1_v_o   (IC_GW_LINK_V    [1])
  ,.p_bsg_link_out1_tkn_i (IC_GW_LINK_TKN  [1])
  ,.p_bsg_link_out1_d0_o  (IC_GW_LINK_D0   [1])
  ,.p_bsg_link_out1_d1_o  (IC_GW_LINK_D1   [1])
  ,.p_bsg_link_out1_d2_o  (IC_GW_LINK_D2   [1])
  ,.p_bsg_link_out1_d3_o  (IC_GW_LINK_D3   [1])
  ,.p_bsg_link_out1_d4_o  (IC_GW_LINK_D4   [1])
  ,.p_bsg_link_out1_d5_o  (IC_GW_LINK_D5   [1])
  ,.p_bsg_link_out1_d6_o  (IC_GW_LINK_D6   [1])
  ,.p_bsg_link_out1_d7_o  (IC_GW_LINK_D7   [1])
  ,.p_bsg_link_out1_d8_o  (IC_GW_LINK_D8   [1])
                          
  ,.p_bsg_link_out2_clk_o (IC_GW_LINK_CLK  [2])
  ,.p_bsg_link_out2_v_o   (IC_GW_LINK_V    [2])
  ,.p_bsg_link_out2_tkn_i (IC_GW_LINK_TKN  [2])
  ,.p_bsg_link_out2_d0_o  (IC_GW_LINK_D0   [2])
  ,.p_bsg_link_out2_d1_o  (IC_GW_LINK_D1   [2])
  ,.p_bsg_link_out2_d2_o  (IC_GW_LINK_D2   [2])
  ,.p_bsg_link_out2_d3_o  (IC_GW_LINK_D3   [2])
  ,.p_bsg_link_out2_d4_o  (IC_GW_LINK_D4   [2])
  ,.p_bsg_link_out2_d5_o  (IC_GW_LINK_D5   [2])
  ,.p_bsg_link_out2_d6_o  (IC_GW_LINK_D6   [2])
  ,.p_bsg_link_out2_d7_o  (IC_GW_LINK_D7   [2])
  ,.p_bsg_link_out2_d8_o  (IC_GW_LINK_D8   [2])
                          
  ,.p_bsg_link_out3_clk_o (IC_GW_LINK_CLK  [3])
  ,.p_bsg_link_out3_v_o   (IC_GW_LINK_V    [3])
  ,.p_bsg_link_out3_tkn_i (IC_GW_LINK_TKN  [3])
  ,.p_bsg_link_out3_d0_o  (IC_GW_LINK_D0   [3])
  ,.p_bsg_link_out3_d1_o  (IC_GW_LINK_D1   [3])
  ,.p_bsg_link_out3_d2_o  (IC_GW_LINK_D2   [3])
  ,.p_bsg_link_out3_d3_o  (IC_GW_LINK_D3   [3])
  ,.p_bsg_link_out3_d4_o  (IC_GW_LINK_D4   [3])
  ,.p_bsg_link_out3_d5_o  (IC_GW_LINK_D5   [3])
  ,.p_bsg_link_out3_d6_o  (IC_GW_LINK_D6   [3])
  ,.p_bsg_link_out3_d7_o  (IC_GW_LINK_D7   [3])
  ,.p_bsg_link_out3_d8_o  (IC_GW_LINK_D8   [3])
                          
  ,.p_bsg_link_out4_clk_o (IC_GW_LINK_CLK  [4])
  ,.p_bsg_link_out4_v_o   (IC_GW_LINK_V    [4])
  ,.p_bsg_link_out4_tkn_i (IC_GW_LINK_TKN  [4])
  ,.p_bsg_link_out4_d0_o  (IC_GW_LINK_D0   [4])
  ,.p_bsg_link_out4_d1_o  (IC_GW_LINK_D1   [4])
  ,.p_bsg_link_out4_d2_o  (IC_GW_LINK_D2   [4])
  ,.p_bsg_link_out4_d3_o  (IC_GW_LINK_D3   [4])
  ,.p_bsg_link_out4_d4_o  (IC_GW_LINK_D4   [4])
  ,.p_bsg_link_out4_d5_o  (IC_GW_LINK_D5   [4])
  ,.p_bsg_link_out4_d6_o  (IC_GW_LINK_D6   [4])
  ,.p_bsg_link_out4_d7_o  (IC_GW_LINK_D7   [4])
  ,.p_bsg_link_out4_d8_o  (IC_GW_LINK_D8   [4])
                          
  ,.p_bsg_link_out5_clk_o (IC_GW_LINK_CLK  [5])
  ,.p_bsg_link_out5_v_o   (IC_GW_LINK_V    [5])
  ,.p_bsg_link_out5_tkn_i (IC_GW_LINK_TKN  [5])
  ,.p_bsg_link_out5_d0_o  (IC_GW_LINK_D0   [5])
  ,.p_bsg_link_out5_d1_o  (IC_GW_LINK_D1   [5])
  ,.p_bsg_link_out5_d2_o  (IC_GW_LINK_D2   [5])
  ,.p_bsg_link_out5_d3_o  (IC_GW_LINK_D3   [5])
  ,.p_bsg_link_out5_d4_o  (IC_GW_LINK_D4   [5])
  ,.p_bsg_link_out5_d5_o  (IC_GW_LINK_D5   [5])
  ,.p_bsg_link_out5_d6_o  (IC_GW_LINK_D6   [5])
  ,.p_bsg_link_out5_d7_o  (IC_GW_LINK_D7   [5])
  ,.p_bsg_link_out5_d8_o  (IC_GW_LINK_D8   [5])
                           
  ,.p_bsg_link_out6_clk_o (IC_GW_LINK_CLK  [6])
  ,.p_bsg_link_out6_v_o   (IC_GW_LINK_V    [6])
  ,.p_bsg_link_out6_tkn_i (IC_GW_LINK_TKN  [6])
  ,.p_bsg_link_out6_d0_o  (IC_GW_LINK_D0   [6])
  ,.p_bsg_link_out6_d1_o  (IC_GW_LINK_D1   [6])
  ,.p_bsg_link_out6_d2_o  (IC_GW_LINK_D2   [6])
  ,.p_bsg_link_out6_d3_o  (IC_GW_LINK_D3   [6])
  ,.p_bsg_link_out6_d4_o  (IC_GW_LINK_D4   [6])
  ,.p_bsg_link_out6_d5_o  (IC_GW_LINK_D5   [6])
  ,.p_bsg_link_out6_d6_o  (IC_GW_LINK_D6   [6])
  ,.p_bsg_link_out6_d7_o  (IC_GW_LINK_D7   [6])
  ,.p_bsg_link_out6_d8_o  (IC_GW_LINK_D8   [6])
                           
  ,.p_bsg_link_out7_clk_o (IC_GW_LINK_CLK  [7])
  ,.p_bsg_link_out7_v_o   (IC_GW_LINK_V    [7])
  ,.p_bsg_link_out7_tkn_i (IC_GW_LINK_TKN  [7])
  ,.p_bsg_link_out7_d0_o  (IC_GW_LINK_D0   [7])
  ,.p_bsg_link_out7_d1_o  (IC_GW_LINK_D1   [7])
  ,.p_bsg_link_out7_d2_o  (IC_GW_LINK_D2   [7])
  ,.p_bsg_link_out7_d3_o  (IC_GW_LINK_D3   [7])
  ,.p_bsg_link_out7_d4_o  (IC_GW_LINK_D4   [7])
  ,.p_bsg_link_out7_d5_o  (IC_GW_LINK_D5   [7])
  ,.p_bsg_link_out7_d6_o  (IC_GW_LINK_D6   [7])
  ,.p_bsg_link_out7_d7_o  (IC_GW_LINK_D7   [7])
  ,.p_bsg_link_out7_d8_o  (IC_GW_LINK_D8   [7])
                           
  ,.p_bsg_link_out8_clk_o (IC_GW_LINK_CLK  [8])
  ,.p_bsg_link_out8_v_o   (IC_GW_LINK_V    [8])
  ,.p_bsg_link_out8_tkn_i (IC_GW_LINK_TKN  [8])
  ,.p_bsg_link_out8_d0_o  (IC_GW_LINK_D0   [8])
  ,.p_bsg_link_out8_d1_o  (IC_GW_LINK_D1   [8])
  ,.p_bsg_link_out8_d2_o  (IC_GW_LINK_D2   [8])
  ,.p_bsg_link_out8_d3_o  (IC_GW_LINK_D3   [8])
  ,.p_bsg_link_out8_d4_o  (IC_GW_LINK_D4   [8])
  ,.p_bsg_link_out8_d5_o  (IC_GW_LINK_D5   [8])
  ,.p_bsg_link_out8_d6_o  (IC_GW_LINK_D6   [8])
  ,.p_bsg_link_out8_d7_o  (IC_GW_LINK_D7   [8])
  ,.p_bsg_link_out8_d8_o  (IC_GW_LINK_D8   [8])
                           
  ,.p_bsg_link_out9_clk_o (IC_GW_LINK_CLK  [9])
  ,.p_bsg_link_out9_v_o   (IC_GW_LINK_V    [9])
  ,.p_bsg_link_out9_tkn_i (IC_GW_LINK_TKN  [9])
  ,.p_bsg_link_out9_d0_o  (IC_GW_LINK_D0   [9])
  ,.p_bsg_link_out9_d1_o  (IC_GW_LINK_D1   [9])
  ,.p_bsg_link_out9_d2_o  (IC_GW_LINK_D2   [9])
  ,.p_bsg_link_out9_d3_o  (IC_GW_LINK_D3   [9])
  ,.p_bsg_link_out9_d4_o  (IC_GW_LINK_D4   [9])
  ,.p_bsg_link_out9_d5_o  (IC_GW_LINK_D5   [9])
  ,.p_bsg_link_out9_d6_o  (IC_GW_LINK_D6   [9])
  ,.p_bsg_link_out9_d7_o  (IC_GW_LINK_D7   [9])
  ,.p_bsg_link_out9_d8_o  (IC_GW_LINK_D8   [9])
                          
  ,.p_bsg_link_out10_clk_o(IC_GW_LINK_CLK  [10])
  ,.p_bsg_link_out10_v_o  (IC_GW_LINK_V    [10])
  ,.p_bsg_link_out10_tkn_i(IC_GW_LINK_TKN  [10])
  ,.p_bsg_link_out10_d0_o (IC_GW_LINK_D0   [10])
  ,.p_bsg_link_out10_d1_o (IC_GW_LINK_D1   [10])
  ,.p_bsg_link_out10_d2_o (IC_GW_LINK_D2   [10])
  ,.p_bsg_link_out10_d3_o (IC_GW_LINK_D3   [10])
  ,.p_bsg_link_out10_d4_o (IC_GW_LINK_D4   [10])
  ,.p_bsg_link_out10_d5_o (IC_GW_LINK_D5   [10])
  ,.p_bsg_link_out10_d6_o (IC_GW_LINK_D6   [10])
  ,.p_bsg_link_out10_d7_o (IC_GW_LINK_D7   [10])
  ,.p_bsg_link_out10_d8_o (IC_GW_LINK_D8   [10])
                           
  ,.p_bsg_link_out11_clk_o(IC_GW_LINK_CLK  [11])
  ,.p_bsg_link_out11_v_o  (IC_GW_LINK_V    [11])
  ,.p_bsg_link_out11_tkn_i(IC_GW_LINK_TKN  [11])
  ,.p_bsg_link_out11_d0_o (IC_GW_LINK_D0   [11])
  ,.p_bsg_link_out11_d1_o (IC_GW_LINK_D1   [11])
  ,.p_bsg_link_out11_d2_o (IC_GW_LINK_D2   [11])
  ,.p_bsg_link_out11_d3_o (IC_GW_LINK_D3   [11])
  ,.p_bsg_link_out11_d4_o (IC_GW_LINK_D4   [11])
  ,.p_bsg_link_out11_d5_o (IC_GW_LINK_D5   [11])
  ,.p_bsg_link_out11_d6_o (IC_GW_LINK_D6   [11])
  ,.p_bsg_link_out11_d7_o (IC_GW_LINK_D7   [11])
  ,.p_bsg_link_out11_d8_o (IC_GW_LINK_D8   [11])
                           
  ,.p_bsg_link_out12_clk_o(IC_GW_LINK_CLK  [12])
  ,.p_bsg_link_out12_v_o  (IC_GW_LINK_V    [12])
  ,.p_bsg_link_out12_tkn_i(IC_GW_LINK_TKN  [12])
  ,.p_bsg_link_out12_d0_o (IC_GW_LINK_D0   [12])
  ,.p_bsg_link_out12_d1_o (IC_GW_LINK_D1   [12])
  ,.p_bsg_link_out12_d2_o (IC_GW_LINK_D2   [12])
  ,.p_bsg_link_out12_d3_o (IC_GW_LINK_D3   [12])
  ,.p_bsg_link_out12_d4_o (IC_GW_LINK_D4   [12])
  ,.p_bsg_link_out12_d5_o (IC_GW_LINK_D5   [12])
  ,.p_bsg_link_out12_d6_o (IC_GW_LINK_D6   [12])
  ,.p_bsg_link_out12_d7_o (IC_GW_LINK_D7   [12])
  ,.p_bsg_link_out12_d8_o (IC_GW_LINK_D8   [12])
                           
  ,.p_bsg_link_out13_clk_o(IC_GW_LINK_CLK  [13])
  ,.p_bsg_link_out13_v_o  (IC_GW_LINK_V    [13])
  ,.p_bsg_link_out13_tkn_i(IC_GW_LINK_TKN  [13])
  ,.p_bsg_link_out13_d0_o (IC_GW_LINK_D0   [13])
  ,.p_bsg_link_out13_d1_o (IC_GW_LINK_D1   [13])
  ,.p_bsg_link_out13_d2_o (IC_GW_LINK_D2   [13])
  ,.p_bsg_link_out13_d3_o (IC_GW_LINK_D3   [13])
  ,.p_bsg_link_out13_d4_o (IC_GW_LINK_D4   [13])
  ,.p_bsg_link_out13_d5_o (IC_GW_LINK_D5   [13])
  ,.p_bsg_link_out13_d6_o (IC_GW_LINK_D6   [13])
  ,.p_bsg_link_out13_d7_o (IC_GW_LINK_D7   [13])
  ,.p_bsg_link_out13_d8_o (IC_GW_LINK_D8   [13])
                           
  ,.p_bsg_link_out14_clk_o(IC_GW_LINK_CLK  [14])
  ,.p_bsg_link_out14_v_o  (IC_GW_LINK_V    [14])
  ,.p_bsg_link_out14_tkn_i(IC_GW_LINK_TKN  [14])
  ,.p_bsg_link_out14_d0_o (IC_GW_LINK_D0   [14])
  ,.p_bsg_link_out14_d1_o (IC_GW_LINK_D1   [14])
  ,.p_bsg_link_out14_d2_o (IC_GW_LINK_D2   [14])
  ,.p_bsg_link_out14_d3_o (IC_GW_LINK_D3   [14])
  ,.p_bsg_link_out14_d4_o (IC_GW_LINK_D4   [14])
  ,.p_bsg_link_out14_d5_o (IC_GW_LINK_D5   [14])
  ,.p_bsg_link_out14_d6_o (IC_GW_LINK_D6   [14])
  ,.p_bsg_link_out14_d7_o (IC_GW_LINK_D7   [14])
  ,.p_bsg_link_out14_d8_o (IC_GW_LINK_D8   [14])
                          
  ,.p_bsg_link_out15_clk_o(IC_GW_LINK_CLK  [15])
  ,.p_bsg_link_out15_v_o  (IC_GW_LINK_V    [15])
  ,.p_bsg_link_out15_tkn_i(IC_GW_LINK_TKN  [15])
  ,.p_bsg_link_out15_d0_o (IC_GW_LINK_D0   [15])
  ,.p_bsg_link_out15_d1_o (IC_GW_LINK_D1   [15])
  ,.p_bsg_link_out15_d2_o (IC_GW_LINK_D2   [15])
  ,.p_bsg_link_out15_d3_o (IC_GW_LINK_D3   [15])
  ,.p_bsg_link_out15_d4_o (IC_GW_LINK_D4   [15])
  ,.p_bsg_link_out15_d5_o (IC_GW_LINK_D5   [15])
  ,.p_bsg_link_out15_d6_o (IC_GW_LINK_D6   [15])
  ,.p_bsg_link_out15_d7_o (IC_GW_LINK_D7   [15])
  ,.p_bsg_link_out15_d8_o (IC_GW_LINK_D8   [15])
                           
  ,.p_bsg_link_out16_clk_o(IC_GW_LINK_CLK  [16])
  ,.p_bsg_link_out16_v_o  (IC_GW_LINK_V    [16])
  ,.p_bsg_link_out16_tkn_i(IC_GW_LINK_TKN  [16])
  ,.p_bsg_link_out16_d0_o (IC_GW_LINK_D0   [16])
  ,.p_bsg_link_out16_d1_o (IC_GW_LINK_D1   [16])
  ,.p_bsg_link_out16_d2_o (IC_GW_LINK_D2   [16])
  ,.p_bsg_link_out16_d3_o (IC_GW_LINK_D3   [16])
  ,.p_bsg_link_out16_d4_o (IC_GW_LINK_D4   [16])
  ,.p_bsg_link_out16_d5_o (IC_GW_LINK_D5   [16])
  ,.p_bsg_link_out16_d6_o (IC_GW_LINK_D6   [16])
  ,.p_bsg_link_out16_d7_o (IC_GW_LINK_D7   [16])
  ,.p_bsg_link_out16_d8_o (IC_GW_LINK_D8   [16])
                           
  ,.p_bsg_link_out17_clk_o(IC_GW_LINK_CLK  [17])
  ,.p_bsg_link_out17_v_o  (IC_GW_LINK_V    [17])
  ,.p_bsg_link_out17_tkn_i(IC_GW_LINK_TKN  [17])
  ,.p_bsg_link_out17_d0_o (IC_GW_LINK_D0   [17])
  ,.p_bsg_link_out17_d1_o (IC_GW_LINK_D1   [17])
  ,.p_bsg_link_out17_d2_o (IC_GW_LINK_D2   [17])
  ,.p_bsg_link_out17_d3_o (IC_GW_LINK_D3   [17])
  ,.p_bsg_link_out17_d4_o (IC_GW_LINK_D4   [17])
  ,.p_bsg_link_out17_d5_o (IC_GW_LINK_D5   [17])
  ,.p_bsg_link_out17_d6_o (IC_GW_LINK_D6   [17])
  ,.p_bsg_link_out17_d7_o (IC_GW_LINK_D7   [17])
  ,.p_bsg_link_out17_d8_o (IC_GW_LINK_D8   [17])
                           
  ,.p_bsg_link_out18_clk_o(IC_GW_LINK_CLK  [18])
  ,.p_bsg_link_out18_v_o  (IC_GW_LINK_V    [18])
  ,.p_bsg_link_out18_tkn_i(IC_GW_LINK_TKN  [18])
  ,.p_bsg_link_out18_d0_o (IC_GW_LINK_D0   [18])
  ,.p_bsg_link_out18_d1_o (IC_GW_LINK_D1   [18])
  ,.p_bsg_link_out18_d2_o (IC_GW_LINK_D2   [18])
  ,.p_bsg_link_out18_d3_o (IC_GW_LINK_D3   [18])
  ,.p_bsg_link_out18_d4_o (IC_GW_LINK_D4   [18])
  ,.p_bsg_link_out18_d5_o (IC_GW_LINK_D5   [18])
  ,.p_bsg_link_out18_d6_o (IC_GW_LINK_D6   [18])
  ,.p_bsg_link_out18_d7_o (IC_GW_LINK_D7   [18])
  ,.p_bsg_link_out18_d8_o (IC_GW_LINK_D8   [18])
                           
  ,.p_bsg_link_out19_clk_o(IC_GW_LINK_CLK  [19])
  ,.p_bsg_link_out19_v_o  (IC_GW_LINK_V    [19])
  ,.p_bsg_link_out19_tkn_i(IC_GW_LINK_TKN  [19])
  ,.p_bsg_link_out19_d0_o (IC_GW_LINK_D0   [19])
  ,.p_bsg_link_out19_d1_o (IC_GW_LINK_D1   [19])
  ,.p_bsg_link_out19_d2_o (IC_GW_LINK_D2   [19])
  ,.p_bsg_link_out19_d3_o (IC_GW_LINK_D3   [19])
  ,.p_bsg_link_out19_d4_o (IC_GW_LINK_D4   [19])
  ,.p_bsg_link_out19_d5_o (IC_GW_LINK_D5   [19])
  ,.p_bsg_link_out19_d6_o (IC_GW_LINK_D6   [19])
  ,.p_bsg_link_out19_d7_o (IC_GW_LINK_D7   [19])
  ,.p_bsg_link_out19_d8_o (IC_GW_LINK_D8   [19])

  ,.p_bsg_tag_clk_i       (GW_TAG_CLKO)
  ,.p_bsg_tag_en_i        (GW_TAG_EN)
  ,.p_bsg_tag_data_i      (GW_TAG_DATAO)
  ,.p_bsg_tag_clk_o       ()
  ,.p_bsg_tag_data_o      ()

  ,.p_clk_A_i             (GW_CLKA)
  ,.p_clk_B_i             (GW_CLKB)
  ,.p_clk_C_i             (GW_CLKC)

  ,.p_clk_o               (IC_CLKO)

  ,.p_sel_0_i             (GW_SEL0)
  ,.p_sel_1_i             (GW_SEL1)
  ,.p_sel_2_i             (GW_SEL2)

  ,.p_clk_async_reset_i   (GW_CLK_RESET)
  ,.p_core_async_reset_i  (GW_CORE_RESET)

  ,.p_misc_o              ()
  );

endmodule
