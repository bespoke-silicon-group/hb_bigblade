module bsg_chip_block (
  output  pad_DL5_0_o_int,      output  pad_DL5_1_o_int,      input   pad_DL5_0_i_int,      input   pad_DL5_1_i_int,
  output  pad_DL5_3_o_int,      output  pad_DL5_2_o_int,      input   pad_DL5_2_i_int,      output  pad_DL5_4_o_int,
  output  pad_DL5_5_o_int,      input   pad_DL5_3_i_int,      input   pad_DL5_4_i_int,      output  pad_DL5_7_o_int,
  output  pad_DL5_6_o_int,      input   pad_DL5_6_i_int,      input   pad_DL5_5_i_int,      output  pad_DL5_9_o_int,
  output  pad_DL5_8_o_int,      input   pad_DL5_7_i_int,      input   pad_DL5_8_i_int,      output  pad_DL5_tkn_o_int,
  output  pad_DL5_10_o_int,     input   pad_DL5_9_i_int,      output  pad_DL5_clk_o_int,    input   pad_DL5_clk_i_int,
  input   pad_DL5_tkn_i_int,    output  pad_DL5_v_o_int,      output  pad_DL5_11_o_int,     input   pad_DL5_v_i_int,
  input   pad_DL5_extra_i_int,  output  pad_DL5_12_o_int,     input   pad_DL5_12_i_int,     input   pad_DL5_11_i_int,
  input   pad_DL5_10_i_int,     output  pad_DL5_13_o_int,     output  pad_DL5_14_o_int,     input   pad_DL5_13_i_int,
  input   pad_DL5_14_i_int,     output  pad_DL5_15_o_int,     output  pad_DL5_extra_o_int,  input   pad_DL5_15_i_int,
  output  pad_DL4_0_o_int,      output  pad_DL4_1_o_int,      input   pad_DL4_0_i_int,      input   pad_DL4_1_i_int,
  output  pad_DL4_3_o_int,      output  pad_DL4_2_o_int,      input   pad_DL4_2_i_int,      output  pad_DL4_4_o_int,
  output  pad_DL4_5_o_int,      input   pad_DL4_3_i_int,      input   pad_DL4_4_i_int,      output  pad_DL4_7_o_int,
  output  pad_DL4_6_o_int,      input   pad_DL4_6_i_int,      input   pad_DL4_5_i_int,      output  pad_DL4_9_o_int,
  output  pad_DL4_8_o_int,      input   pad_DL4_7_i_int,      input   pad_DL4_8_i_int,      output  pad_DL4_tkn_o_int,
  output  pad_DL4_10_o_int,     input   pad_DL4_9_i_int,      output  pad_DL4_clk_o_int,    input   pad_DL4_clk_i_int,
  input   pad_DL4_tkn_i_int,    output  pad_DL4_v_o_int,      output  pad_DL4_11_o_int,     input   pad_DL4_v_i_int,
  input   pad_DL4_extra_i_int,  output  pad_DL4_12_o_int,     input   pad_DL4_12_i_int,     input   pad_DL4_11_i_int,
  input   pad_DL4_10_i_int,     output  pad_DL4_13_o_int,     output  pad_DL4_14_o_int,     input   pad_DL4_13_i_int,
  input   pad_DL4_14_i_int,     output  pad_DL4_15_o_int,     output  pad_DL4_extra_o_int,  input   pad_DL4_15_i_int,
  output  pad_DL3_0_o_int,      output  pad_DL3_1_o_int,      input   pad_DL3_0_i_int,      input   pad_DL3_1_i_int,
  output  pad_DL3_3_o_int,      output  pad_DL3_2_o_int,      input   pad_DL3_2_i_int,      output  pad_DL3_4_o_int,
  output  pad_DL3_5_o_int,      input   pad_DL3_3_i_int,      input   pad_DL3_4_i_int,      output  pad_DL3_7_o_int,
  output  pad_DL3_6_o_int,      input   pad_DL3_6_i_int,      input   pad_DL3_5_i_int,      output  pad_DL3_9_o_int,
  output  pad_DL3_8_o_int,      input   pad_DL3_7_i_int,      input   pad_DL3_8_i_int,      output  pad_DL3_tkn_o_int,
  output  pad_DL3_10_o_int,     input   pad_DL3_9_i_int,      output  pad_DL3_clk_o_int,    input   pad_DL3_clk_i_int,
  input   pad_DL3_tkn_i_int,    output  pad_DL3_v_o_int,      output  pad_DL3_11_o_int,     input   pad_DL3_v_i_int,
  input   pad_DL3_extra_i_int,  output  pad_DL3_12_o_int,     input   pad_DL3_12_i_int,     input   pad_DL3_11_i_int,
  input   pad_DL3_10_i_int,     output  pad_DL3_13_o_int,     output  pad_DL3_14_o_int,     input   pad_DL3_13_i_int,
  input   pad_DL3_14_i_int,     output  pad_DL3_15_o_int,     output  pad_DL3_extra_o_int,  input   pad_DL3_15_i_int,
  output  pad_DL2_0_o_int,      output  pad_DL2_1_o_int,      input   pad_DL2_0_i_int,      input   pad_DL2_1_i_int,
  output  pad_DL2_3_o_int,      output  pad_DL2_2_o_int,      input   pad_DL2_2_i_int,      output  pad_DL2_4_o_int,
  output  pad_DL2_5_o_int,      input   pad_DL2_3_i_int,      input   pad_DL2_4_i_int,      output  pad_DL2_7_o_int,
  output  pad_DL2_6_o_int,      input   pad_DL2_6_i_int,      input   pad_DL2_5_i_int,      output  pad_DL2_9_o_int,
  output  pad_DL2_8_o_int,      input   pad_DL2_7_i_int,      input   pad_DL2_8_i_int,      output  pad_DL2_tkn_o_int,
  output  pad_DL2_10_o_int,     input   pad_DL2_9_i_int,      output  pad_DL2_clk_o_int,    input   pad_DL2_clk_i_int,
  input   pad_DL2_tkn_i_int,    output  pad_DL2_v_o_int,      output  pad_DL2_11_o_int,     input   pad_DL2_v_i_int,
  input   pad_DL2_extra_i_int,  output  pad_DL2_12_o_int,     input   pad_DL2_12_i_int,     input   pad_DL2_11_i_int,
  input   pad_DL2_10_i_int,     output  pad_DL2_13_o_int,     output  pad_DL2_14_o_int,     input   pad_DL2_13_i_int,
  input   pad_DL2_14_i_int,     output  pad_DL2_15_o_int,     output  pad_DL2_extra_o_int,  input   pad_DL2_15_i_int,
  output  pad_DL1_0_o_int,      output  pad_DL1_1_o_int,      input   pad_DL1_0_i_int,      input   pad_DL1_1_i_int,
  output  pad_DL1_3_o_int,      output  pad_DL1_2_o_int,      input   pad_DL1_2_i_int,      output  pad_DL1_4_o_int,
  output  pad_DL1_5_o_int,      input   pad_DL1_3_i_int,      input   pad_DL1_4_i_int,      output  pad_DL1_7_o_int,
  output  pad_DL1_6_o_int,      input   pad_DL1_6_i_int,      input   pad_DL1_5_i_int,      output  pad_DL1_9_o_int,
  output  pad_DL1_8_o_int,      input   pad_DL1_7_i_int,      input   pad_DL1_8_i_int,      output  pad_DL1_tkn_o_int,
  output  pad_DL1_10_o_int,     input   pad_DL1_9_i_int,      output  pad_DL1_clk_o_int,    input   pad_DL1_clk_i_int,
  input   pad_DL1_tkn_i_int,    output  pad_DL1_v_o_int,      output  pad_DL1_11_o_int,     input   pad_DL1_v_i_int,
  input   pad_DL1_extra_i_int,  output  pad_DL1_12_o_int,     input   pad_DL1_12_i_int,     input   pad_DL1_11_i_int,
  input   pad_DL1_10_i_int,     output  pad_DL1_13_o_int,     output  pad_DL1_14_o_int,     input   pad_DL1_13_i_int,
  input   pad_DL1_14_i_int,     output  pad_DL1_15_o_int,     output  pad_DL1_extra_o_int,  input   pad_DL1_15_i_int,
  input   pad_ML0_0_i_int,      input   pad_ML0_1_i_int,      input   pad_ML0_2_i_int,      input   pad_ML0_6_i_int,
  input   pad_ML0_5_i_int,      input   pad_ML0_3_i_int,      input   pad_ML0_4_i_int,      output  pad_DL0_0_o_int,
  output  pad_DL0_1_o_int,      input   pad_DL0_0_i_int,      input   pad_DL0_1_i_int,      output  pad_DL0_3_o_int,
  output  pad_DL0_2_o_int,      input   pad_DL0_2_i_int,      output  pad_DL0_4_o_int,      output  pad_DL0_5_o_int,
  input   pad_DL0_3_i_int,      input   pad_DL0_4_i_int,      output  pad_DL0_7_o_int,      output  pad_DL0_6_o_int,
  input   pad_DL0_6_i_int,      input   pad_DL0_5_i_int,      output  pad_DL0_9_o_int,      output  pad_DL0_8_o_int,
  input   pad_DL0_7_i_int,      input   pad_DL0_8_i_int,      output  pad_DL0_tkn_o_int,    output  pad_DL0_10_o_int,
  input   pad_DL0_9_i_int,      output  pad_DL0_clk_o_int,    input   pad_DL0_clk_i_int,    input   pad_DL0_tkn_i_int,
  output  pad_DL0_v_o_int,      output  pad_DL0_11_o_int,     input   pad_DL0_v_i_int,      input   pad_DL0_extra_i_int,
  output  pad_DL0_12_o_int,     input   pad_DL0_12_i_int,     input   pad_DL0_11_i_int,     input   pad_DL0_10_i_int,
  output  pad_DL0_13_o_int,     output  pad_DL0_14_o_int,     input   pad_DL0_13_i_int,     input   pad_DL0_14_i_int,
  output  pad_DL0_15_o_int,     output  pad_DL0_extra_o_int,  input   pad_DL0_15_i_int,     output  pad_IT0_0_o_int,
  output  pad_IT0_1_o_int,      input   pad_IT0_0_i_int,      input   pad_IT0_1_i_int,      output  pad_IT0_3_o_int,
  output  pad_IT0_2_o_int,      input   pad_IT0_2_i_int,      output  pad_IT0_4_o_int,      output  pad_IT0_5_o_int,
  input   pad_IT0_3_i_int,      input   pad_IT0_4_i_int,      output  pad_IT0_7_o_int,      output  pad_IT0_6_o_int,
  input   pad_IT0_6_i_int,      input   pad_IT0_5_i_int,      output  pad_IT0_9_o_int,      output  pad_IT0_8_o_int,
  input   pad_IT0_7_i_int,      input   pad_IT0_8_i_int,      output  pad_IT0_tkn_o_int,    output  pad_IT0_10_o_int,
  input   pad_IT0_9_i_int,      output  pad_IT0_clk_o_int,    input   pad_IT0_clk_i_int,    input   pad_IT0_tkn_i_int,
  output  pad_IT0_v_o_int,      output  pad_IT0_11_o_int,     input   pad_IT0_v_i_int,      input   pad_IT0_extra_i_int,
  output  pad_IT0_12_o_int,     input   pad_IT0_12_i_int,     input   pad_IT0_11_i_int,     input   pad_IT0_10_i_int,
  output  pad_IT0_13_o_int,     output  pad_IT0_14_o_int,     input   pad_IT0_13_i_int,     input   pad_IT0_14_i_int,
  output  pad_IT0_15_o_int,     output  pad_IT0_extra_o_int,  input   pad_IT0_15_i_int,     output  pad_CT0_0_o_int,
  output  pad_CT0_1_o_int,      input   pad_CT0_0_i_int,      input   pad_CT0_1_i_int,      output  pad_CT0_2_o_int,
  output  pad_CT0_tkn_o_int,    input   pad_CT0_2_i_int,      output  pad_CT0_clk_o_int,    output  pad_CT0_3_o_int,
  input   pad_CT0_clk_i_int,    input   pad_CT0_3_i_int,      output  pad_CT0_4_o_int,      input   pad_CT0_v_i_int,
  input   pad_CT0_4_i_int,      input   pad_CT0_tkn_i_int,    output  pad_CT0_5_o_int,      output  pad_CT0_6_o_int,
  input   pad_CT0_5_i_int,      input   pad_CT0_6_i_int,      output  pad_CT0_7_o_int,      output  pad_CT0_v_o_int,
  input   pad_CT0_7_i_int,      output  pad_IT1_0_o_int,      output  pad_IT1_1_o_int,      input   pad_IT1_0_i_int,
  input   pad_IT1_1_i_int,      output  pad_IT1_3_o_int,      output  pad_IT1_2_o_int,      input   pad_IT1_2_i_int,
  output  pad_IT1_4_o_int,      output  pad_IT1_5_o_int,      input   pad_IT1_3_i_int,      input   pad_IT1_4_i_int,
  output  pad_IT1_7_o_int,      output  pad_IT1_6_o_int,      input   pad_IT1_6_i_int,      input   pad_IT1_5_i_int,
  output  pad_IT1_9_o_int,      output  pad_IT1_8_o_int,      input   pad_IT1_7_i_int,      input   pad_IT1_8_i_int,
  output  pad_IT1_tkn_o_int,    output  pad_IT1_10_o_int,     input   pad_IT1_9_i_int,      output  pad_IT1_clk_o_int,
  input   pad_IT1_clk_i_int,    input   pad_IT1_tkn_i_int,    output  pad_IT1_v_o_int,      output  pad_IT1_11_o_int,
  input   pad_IT1_v_i_int,      input   pad_IT1_extra_i_int,  output  pad_IT1_12_o_int,     input   pad_IT1_12_i_int,
  input   pad_IT1_11_i_int,     input   pad_IT1_10_i_int,     output  pad_IT1_13_o_int,     output  pad_IT1_14_o_int,
  input   pad_IT1_13_i_int,     input   pad_IT1_14_i_int,     output  pad_IT1_15_o_int,     output  pad_IT1_extra_o_int,
  input   pad_IT1_15_i_int,     output  pad_DR0_0_o_int,      output  pad_DR0_1_o_int,      input   pad_DR0_0_i_int,
  input   pad_DR0_1_i_int,      output  pad_DR0_3_o_int,      output  pad_DR0_2_o_int,      input   pad_DR0_2_i_int,
  output  pad_DR0_4_o_int,      output  pad_DR0_5_o_int,      input   pad_DR0_3_i_int,      input   pad_DR0_4_i_int,
  output  pad_DR0_7_o_int,      output  pad_DR0_6_o_int,      input   pad_DR0_6_i_int,      input   pad_DR0_5_i_int,
  output  pad_DR0_9_o_int,      output  pad_DR0_8_o_int,      input   pad_DR0_7_i_int,      input   pad_DR0_8_i_int,
  output  pad_DR0_tkn_o_int,    output  pad_DR0_10_o_int,     input   pad_DR0_9_i_int,      output  pad_DR0_clk_o_int,
  input   pad_DR0_clk_i_int,    input   pad_DR0_tkn_i_int,    output  pad_DR0_v_o_int,      output  pad_DR0_11_o_int,
  input   pad_DR0_v_i_int,      input   pad_DR0_extra_i_int,  output  pad_DR0_12_o_int,     input   pad_DR0_12_i_int,
  input   pad_DR0_11_i_int,     input   pad_DR0_10_i_int,     output  pad_DR0_13_o_int,     output  pad_DR0_14_o_int,
  input   pad_DR0_13_i_int,     input   pad_DR0_14_i_int,     output  pad_DR0_15_o_int,     output  pad_DR0_extra_o_int,
  input   pad_DR0_15_i_int,     input   pad_MR0_2_i_int,      input   pad_MR0_1_i_int,      input   pad_MR0_0_i_int,
  input   pad_DR1_15_i_int,     output  pad_DR1_extra_o_int,  output  pad_DR1_15_o_int,     input   pad_DR1_14_i_int,
  input   pad_DR1_13_i_int,     output  pad_DR1_14_o_int,     output  pad_DR1_13_o_int,     input   pad_DR1_10_i_int,
  input   pad_DR1_11_i_int,     input   pad_DR1_12_i_int,     output  pad_DR1_12_o_int,     input   pad_DR1_extra_i_int,
  input   pad_DR1_v_i_int,      output  pad_DR1_11_o_int,     output  pad_DR1_v_o_int,      input   pad_DR1_tkn_i_int,
  input   pad_DR1_clk_i_int,    output  pad_DR1_clk_o_int,    input   pad_DR1_9_i_int,      output  pad_DR1_10_o_int,
  output  pad_DR1_tkn_o_int,    input   pad_DR1_8_i_int,      input   pad_DR1_7_i_int,      output  pad_DR1_8_o_int,
  output  pad_DR1_9_o_int,      input   pad_DR1_5_i_int,      input   pad_DR1_6_i_int,      output  pad_DR1_6_o_int,
  output  pad_DR1_7_o_int,      input   pad_DR1_4_i_int,      input   pad_DR1_3_i_int,      output  pad_DR1_5_o_int,
  output  pad_DR1_4_o_int,      input   pad_DR1_2_i_int,      output  pad_DR1_2_o_int,      output  pad_DR1_3_o_int,
  input   pad_DR1_1_i_int,      input   pad_DR1_0_i_int,      output  pad_DR1_1_o_int,      output  pad_DR1_0_o_int,
  input   pad_DR2_15_i_int,     output  pad_DR2_extra_o_int,  output  pad_DR2_15_o_int,     input   pad_DR2_14_i_int,
  input   pad_DR2_13_i_int,     output  pad_DR2_14_o_int,     output  pad_DR2_13_o_int,     input   pad_DR2_10_i_int,
  input   pad_DR2_11_i_int,     input   pad_DR2_12_i_int,     output  pad_DR2_12_o_int,     input   pad_DR2_extra_i_int,
  input   pad_DR2_v_i_int,      output  pad_DR2_11_o_int,     output  pad_DR2_v_o_int,      input   pad_DR2_tkn_i_int,
  input   pad_DR2_clk_i_int,    output  pad_DR2_clk_o_int,    input   pad_DR2_9_i_int,      output  pad_DR2_10_o_int,
  output  pad_DR2_tkn_o_int,    input   pad_DR2_8_i_int,      input   pad_DR2_7_i_int,      output  pad_DR2_8_o_int,
  output  pad_DR2_9_o_int,      input   pad_DR2_5_i_int,      input   pad_DR2_6_i_int,      output  pad_DR2_6_o_int,
  output  pad_DR2_7_o_int,      input   pad_DR2_4_i_int,      input   pad_DR2_3_i_int,      output  pad_DR2_5_o_int,
  output  pad_DR2_4_o_int,      input   pad_DR2_2_i_int,      output  pad_DR2_2_o_int,      output  pad_DR2_3_o_int,
  input   pad_DR2_1_i_int,      input   pad_DR2_0_i_int,      output  pad_DR2_1_o_int,      output  pad_DR2_0_o_int,
  input   pad_DR3_15_i_int,     output  pad_DR3_extra_o_int,  output  pad_DR3_15_o_int,     input   pad_DR3_14_i_int,
  input   pad_DR3_13_i_int,     output  pad_DR3_14_o_int,     output  pad_DR3_13_o_int,     input   pad_DR3_10_i_int,
  input   pad_DR3_11_i_int,     input   pad_DR3_12_i_int,     output  pad_DR3_12_o_int,     input   pad_DR3_extra_i_int,
  input   pad_DR3_v_i_int,      output  pad_DR3_11_o_int,     output  pad_DR3_v_o_int,      input   pad_DR3_tkn_i_int,
  input   pad_DR3_clk_i_int,    output  pad_DR3_clk_o_int,    input   pad_DR3_9_i_int,      output  pad_DR3_10_o_int,
  output  pad_DR3_tkn_o_int,    input   pad_DR3_8_i_int,      input   pad_DR3_7_i_int,      output  pad_DR3_8_o_int,
  output  pad_DR3_9_o_int,      input   pad_DR3_5_i_int,      input   pad_DR3_6_i_int,      output  pad_DR3_6_o_int,
  output  pad_DR3_7_o_int,      input   pad_DR3_4_i_int,      input   pad_DR3_3_i_int,      output  pad_DR3_5_o_int,
  output  pad_DR3_4_o_int,      input   pad_DR3_2_i_int,      output  pad_DR3_2_o_int,      output  pad_DR3_3_o_int,
  input   pad_DR3_1_i_int,      input   pad_DR3_0_i_int,      output  pad_DR3_1_o_int,      output  pad_DR3_0_o_int,
  input   pad_DR4_15_i_int,     output  pad_DR4_extra_o_int,  output  pad_DR4_15_o_int,     input   pad_DR4_14_i_int,
  input   pad_DR4_13_i_int,     output  pad_DR4_14_o_int,     output  pad_DR4_13_o_int,     input   pad_DR4_10_i_int,
  input   pad_DR4_11_i_int,     input   pad_DR4_12_i_int,     output  pad_DR4_12_o_int,     input   pad_DR4_extra_i_int,
  input   pad_DR4_v_i_int,      output  pad_DR4_11_o_int,     output  pad_DR4_v_o_int,      input   pad_DR4_tkn_i_int,
  input   pad_DR4_clk_i_int,    output  pad_DR4_clk_o_int,    input   pad_DR4_9_i_int,      output  pad_DR4_10_o_int,
  output  pad_DR4_tkn_o_int,    input   pad_DR4_8_i_int,      input   pad_DR4_7_i_int,      output  pad_DR4_8_o_int,
  output  pad_DR4_9_o_int,      input   pad_DR4_5_i_int,      input   pad_DR4_6_i_int,      output  pad_DR4_6_o_int,
  output  pad_DR4_7_o_int,      input   pad_DR4_4_i_int,      input   pad_DR4_3_i_int,      output  pad_DR4_5_o_int,
  output  pad_DR4_4_o_int,      input   pad_DR4_2_i_int,      output  pad_DR4_2_o_int,      output  pad_DR4_3_o_int,
  input   pad_DR4_1_i_int,      input   pad_DR4_0_i_int,      output  pad_DR4_1_o_int,      output  pad_DR4_0_o_int,
  input   pad_DR5_15_i_int,     output  pad_DR5_extra_o_int,  output  pad_DR5_15_o_int,     input   pad_DR5_14_i_int,
  input   pad_DR5_13_i_int,     output  pad_DR5_14_o_int,     output  pad_DR5_13_o_int,     input   pad_DR5_10_i_int,
  input   pad_DR5_11_i_int,     input   pad_DR5_12_i_int,     output  pad_DR5_12_o_int,     input   pad_DR5_extra_i_int,
  input   pad_DR5_v_i_int,      output  pad_DR5_11_o_int,     output  pad_DR5_v_o_int,      input   pad_DR5_tkn_i_int,
  input   pad_DR5_clk_i_int,    output  pad_DR5_clk_o_int,    input   pad_DR5_9_i_int,      output  pad_DR5_10_o_int,
  output  pad_DR5_tkn_o_int,    input   pad_DR5_8_i_int,      input   pad_DR5_7_i_int,      output  pad_DR5_8_o_int,
  output  pad_DR5_9_o_int,      input   pad_DR5_5_i_int,      input   pad_DR5_6_i_int,      output  pad_DR5_6_o_int,
  output  pad_DR5_7_o_int,      input   pad_DR5_4_i_int,      input   pad_DR5_3_i_int,      output  pad_DR5_5_o_int,
  output  pad_DR5_4_o_int,      input   pad_DR5_2_i_int,      output  pad_DR5_2_o_int,      output  pad_DR5_3_o_int,
  input   pad_DR5_1_i_int,      input   pad_DR5_0_i_int,      output  pad_DR5_1_o_int,      output  pad_DR5_0_o_int,
  input   pad_MR1_5_i_int,      input   pad_MR1_6_i_int,      input   pad_MR1_7_i_int,      input   pad_MR1_4_i_int,
  input   pad_MR1_3_i_int,      input   pad_MR1_0_i_int,      input   pad_MR1_1_i_int,      input   pad_MR1_2_i_int,
  input   pad_DR6_15_i_int,     output  pad_DR6_extra_o_int,  output  pad_DR6_15_o_int,     input   pad_DR6_14_i_int,
  input   pad_DR6_13_i_int,     output  pad_DR6_14_o_int,     output  pad_DR6_13_o_int,     input   pad_DR6_10_i_int,
  input   pad_DR6_11_i_int,     input   pad_DR6_12_i_int,     output  pad_DR6_12_o_int,     input   pad_DR6_extra_i_int,
  input   pad_DR6_v_i_int,      output  pad_DR6_11_o_int,     output  pad_DR6_v_o_int,      input   pad_DR6_tkn_i_int,
  input   pad_DR6_clk_i_int,    output  pad_DR6_clk_o_int,    input   pad_DR6_9_i_int,      output  pad_DR6_10_o_int,
  output  pad_DR6_tkn_o_int,    input   pad_DR6_8_i_int,      input   pad_DR6_7_i_int,      output  pad_DR6_8_o_int,
  output  pad_DR6_9_o_int,      input   pad_DR6_5_i_int,      input   pad_DR6_6_i_int,      output  pad_DR6_6_o_int,
  output  pad_DR6_7_o_int,      input   pad_DR6_4_i_int,      input   pad_DR6_3_i_int,      output  pad_DR6_5_o_int,
  output  pad_DR6_4_o_int,      input   pad_DR6_2_i_int,      output  pad_DR6_2_o_int,      output  pad_DR6_3_o_int,
  input   pad_DR6_1_i_int,      input   pad_DR6_0_i_int,      output  pad_DR6_1_o_int,      output  pad_DR6_0_o_int,
  input   pad_DR7_15_i_int,     output  pad_DR7_extra_o_int,  output  pad_DR7_15_o_int,     input   pad_DR7_14_i_int,
  input   pad_DR7_13_i_int,     output  pad_DR7_14_o_int,     output  pad_DR7_13_o_int,     input   pad_DR7_10_i_int,
  input   pad_DR7_11_i_int,     input   pad_DR7_12_i_int,     output  pad_DR7_12_o_int,     input   pad_DR7_extra_i_int,
  input   pad_DR7_v_i_int,      output  pad_DR7_11_o_int,     output  pad_DR7_v_o_int,      input   pad_DR7_tkn_i_int,
  input   pad_DR7_clk_i_int,    output  pad_DR7_clk_o_int,    input   pad_DR7_9_i_int,      output  pad_DR7_10_o_int,
  output  pad_DR7_tkn_o_int,    input   pad_DR7_8_i_int,      input   pad_DR7_7_i_int,      output  pad_DR7_8_o_int,
  output  pad_DR7_9_o_int,      input   pad_DR7_5_i_int,      input   pad_DR7_6_i_int,      output  pad_DR7_6_o_int,
  output  pad_DR7_7_o_int,      input   pad_DR7_4_i_int,      input   pad_DR7_3_i_int,      output  pad_DR7_5_o_int,
  output  pad_DR7_4_o_int,      input   pad_DR7_2_i_int,      output  pad_DR7_2_o_int,      output  pad_DR7_3_o_int,
  input   pad_DR7_1_i_int,      input   pad_DR7_0_i_int,      output  pad_DR7_1_o_int,      output  pad_DR7_0_o_int,
  input   pad_CB0_7_i_int,      output  pad_CB0_v_o_int,      output  pad_CB0_7_o_int,      input   pad_CB0_6_i_int,
  input   pad_CB0_5_i_int,      output  pad_CB0_6_o_int,      output  pad_CB0_5_o_int,      input   pad_CB0_tkn_i_int,
  input   pad_CB0_4_i_int,      input   pad_CB0_v_i_int,      output  pad_CB0_4_o_int,      input   pad_CB0_3_i_int,
  input   pad_CB0_clk_i_int,    output  pad_CB0_3_o_int,      output  pad_CB0_clk_o_int,    input   pad_CB0_2_i_int,
  output  pad_CB0_tkn_o_int,    output  pad_CB0_2_o_int,      input   pad_CB0_1_i_int,      input   pad_CB0_0_i_int,
  output  pad_CB0_1_o_int,      output  pad_CB0_0_o_int,      input   pad_DL7_15_i_int,     output  pad_DL7_extra_o_int,
  output  pad_DL7_15_o_int,     input   pad_DL7_14_i_int,     input   pad_DL7_13_i_int,     output  pad_DL7_14_o_int,
  output  pad_DL7_13_o_int,     input   pad_DL7_10_i_int,     input   pad_DL7_11_i_int,     input   pad_DL7_12_i_int,
  output  pad_DL7_12_o_int,     input   pad_DL7_extra_i_int,  input   pad_DL7_v_i_int,      output  pad_DL7_11_o_int,
  output  pad_DL7_v_o_int,      input   pad_DL7_tkn_i_int,    input   pad_DL7_clk_i_int,    output  pad_DL7_clk_o_int,
  input   pad_DL7_9_i_int,      output  pad_DL7_10_o_int,     output  pad_DL7_tkn_o_int,    input   pad_DL7_8_i_int,
  input   pad_DL7_7_i_int,      output  pad_DL7_8_o_int,      output  pad_DL7_9_o_int,      input   pad_DL7_5_i_int,
  input   pad_DL7_6_i_int,      output  pad_DL7_6_o_int,      output  pad_DL7_7_o_int,      input   pad_DL7_4_i_int,
  input   pad_DL7_3_i_int,      output  pad_DL7_5_o_int,      output  pad_DL7_4_o_int,      input   pad_DL7_2_i_int,
  output  pad_DL7_2_o_int,      output  pad_DL7_3_o_int,      input   pad_DL7_1_i_int,      input   pad_DL7_0_i_int,
  output  pad_DL7_1_o_int,      output  pad_DL7_0_o_int,      input   pad_DL6_15_i_int,     output  pad_DL6_extra_o_int,
  output  pad_DL6_15_o_int,     input   pad_DL6_14_i_int,     input   pad_DL6_13_i_int,     output  pad_DL6_14_o_int,
  output  pad_DL6_13_o_int,     input   pad_DL6_10_i_int,     input   pad_DL6_11_i_int,     input   pad_DL6_12_i_int,
  output  pad_DL6_12_o_int,     input   pad_DL6_extra_i_int,  input   pad_DL6_v_i_int,      output  pad_DL6_11_o_int,
  output  pad_DL6_v_o_int,      input   pad_DL6_tkn_i_int,    input   pad_DL6_clk_i_int,    output  pad_DL6_clk_o_int,
  input   pad_DL6_9_i_int,      output  pad_DL6_10_o_int,     output  pad_DL6_tkn_o_int,    input   pad_DL6_8_i_int,
  input   pad_DL6_7_i_int,      output  pad_DL6_8_o_int,      output  pad_DL6_9_o_int,      input   pad_DL6_5_i_int,
  input   pad_DL6_6_i_int,      output  pad_DL6_6_o_int,      output  pad_DL6_7_o_int,      input   pad_DL6_4_i_int,
  input   pad_DL6_3_i_int,      output  pad_DL6_5_o_int,      output  pad_DL6_4_o_int,      input   pad_DL6_2_i_int,
  output  pad_DL6_2_o_int,      output  pad_DL6_3_o_int,      input   pad_DL6_1_i_int,      input   pad_DL6_0_i_int,
  output  pad_DL6_1_o_int,      output  pad_DL6_0_o_int,      input   pad_ML1_2_i_int,      input   pad_ML1_1_i_int,
  input   pad_ML1_0_i_int
);


endmodule
