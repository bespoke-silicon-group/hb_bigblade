../../bigblade_bp_unicore/v/bp_cce_to_mc_bridge.sv