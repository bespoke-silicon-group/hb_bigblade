module bsg_manycore_link_to_sdr_north
`include "bsg_manycore_link_to_sdr.v"
endmodule