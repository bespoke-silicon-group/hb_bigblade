//
// This is a blackbox for the bsg_chip_block which can be found in the
// bigbalde_toplevel_block design directory.
//

`include "bsg_padmapping.v"
`include "bsg_iopad_macros.v"

module bsg_chip_block

`include "bsg_chip_block_pinout.v"

endmodule
