module bsg_manycore_link_to_sdr_south
`include "bsg_manycore_link_to_sdr.v"
endmodule