 instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow liblist `BSG_MANYCORE_LINK_SDR_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_0__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_1__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_2__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.mc_y_3__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_0__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_0__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_1__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_2__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.mc_y_3__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_1__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_0__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_1__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_2__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.mc_y_3__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_2__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.north_vc_x_0__north_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_0__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_1__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_2__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_0__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;   
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_0__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_1__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_2__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_3__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_4__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_5__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_6__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_7__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_8__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_9__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_10__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_11__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_12__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_13__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_14__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.mc_y_3__mc_x_0__mc.y_1__x_15__tile liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME; 
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_0__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_1__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_2__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_3__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_4__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_5__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_6__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_7__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_8__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_9__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_10__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_11__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_12__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_13__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_14__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;  
instance bsg_bigblade_pcb.IC.ASIC.block.core_complex_core_0__podrow.podrow.px_3__pod.south_vc_x_0__south_vc_row.vc_y_0__vc_x_15__vc liblist `BSG_MANYCORE_TILE_LIBRARY_NAME `BSG_CHIP_LIBRARY_NAME;

